`include "typedef.vh"
/*module sigma_int(input data_type in,
	 output data_type out);
	 	 always_comb
	 	 	 if (in[16:0] >= 0 && in <= 2) out = 2047;
	 	 	 else if (in[16:0] >= 3 && in <= 6) out = 2048;
	 	 	 else if (in[16:0] >= 7 && in <= 10) out = 2049;
	 	 	 else if (in[16:0] >= 11 && in <= 14) out = 2050;
	 	 	 else if (in[16:0] >= 15 && in <= 18) out = 2051;
	 	 	 else if (in[16:0] >= 19 && in <= 22) out = 2052;
	 	 	 else if (in[16:0] >= 23 && in <= 26) out = 2053;
	 	 	 else if (in[16:0] >= 27 && in <= 30) out = 2054;
	 	 	 else if (in[16:0] >= 31 && in <= 34) out = 2055;
	 	 	 else if (in[16:0] >= 35 && in <= 38) out = 2056;
	 	 	 else if (in[16:0] >= 39 && in <= 42) out = 2057;
	 	 	 else if (in[16:0] >= 43 && in <= 46) out = 2058;
	 	 	 else if (in[16:0] >= 47 && in <= 50) out = 2059;
	 	 	 else if (in[16:0] >= 51 && in <= 54) out = 2060;
	 	 	 else if (in[16:0] >= 55 && in <= 58) out = 2061;
	 	 	 else if (in[16:0] >= 59 && in <= 62) out = 2062;
	 	 	 else if (in[16:0] >= 63 && in <= 66) out = 2063;
	 	 	 else if (in[16:0] >= 67 && in <= 70) out = 2064;
	 	 	 else if (in[16:0] >= 71 && in <= 74) out = 2065;
	 	 	 else if (in[16:0] >= 75 && in <= 78) out = 2066;
	 	 	 else if (in[16:0] >= 79 && in <= 82) out = 2067;
	 	 	 else if (in[16:0] >= 83 && in <= 86) out = 2068;
	 	 	 else if (in[16:0] >= 87 && in <= 90) out = 2069;
	 	 	 else if (in[16:0] >= 91 && in <= 94) out = 2070;
	 	 	 else if (in[16:0] >= 95 && in <= 98) out = 2071;
	 	 	 else if (in[16:0] >= 99 && in <= 102) out = 2072;
	 	 	 else if (in[16:0] >= 103 && in <= 106) out = 2073;
	 	 	 else if (in[16:0] >= 107 && in <= 110) out = 2074;
	 	 	 else if (in[16:0] >= 111 && in <= 114) out = 2075;
	 	 	 else if (in[16:0] >= 115 && in <= 118) out = 2076;
	 	 	 else if (in[16:0] >= 119 && in <= 122) out = 2077;
	 	 	 else if (in[16:0] >= 123 && in <= 126) out = 2078;
	 	 	 else if (in[16:0] >= 127 && in <= 130) out = 2079;
	 	 	 else if (in[16:0] >= 131 && in <= 134) out = 2080;
	 	 	 else if (in[16:0] >= 135 && in <= 138) out = 2081;
	 	 	 else if (in[16:0] >= 139 && in <= 142) out = 2082;
	 	 	 else if (in[16:0] >= 143 && in <= 146) out = 2083;
	 	 	 else if (in[16:0] >= 147 && in <= 150) out = 2084;
	 	 	 else if (in[16:0] >= 151 && in <= 154) out = 2085;
	 	 	 else if (in[16:0] >= 155 && in <= 158) out = 2086;
	 	 	 else if (in[16:0] >= 159 && in <= 162) out = 2087;
	 	 	 else if (in[16:0] >= 163 && in <= 166) out = 2088;
	 	 	 else if (in[16:0] >= 167 && in <= 170) out = 2089;
	 	 	 else if (in[16:0] >= 171 && in <= 174) out = 2090;
	 	 	 else if (in[16:0] >= 175 && in <= 178) out = 2091;
	 	 	 else if (in[16:0] >= 179 && in <= 182) out = 2092;
	 	 	 else if (in[16:0] >= 183 && in <= 186) out = 2093;
	 	 	 else if (in[16:0] >= 187 && in <= 190) out = 2094;
	 	 	 else if (in[16:0] >= 191 && in <= 194) out = 2095;
	 	 	 else if (in[16:0] >= 195 && in <= 198) out = 2096;
	 	 	 else if (in[16:0] >= 199 && in <= 202) out = 2097;
	 	 	 else if (in[16:0] >= 203 && in <= 206) out = 2098;
	 	 	 else if (in[16:0] >= 207 && in <= 210) out = 2099;
	 	 	 else if (in[16:0] >= 211 && in <= 214) out = 2100;
	 	 	 else if (in[16:0] >= 215 && in <= 218) out = 2101;
	 	 	 else if (in[16:0] >= 219 && in <= 222) out = 2102;
	 	 	 else if (in[16:0] >= 223 && in <= 226) out = 2103;
	 	 	 else if (in[16:0] >= 227 && in <= 230) out = 2104;
	 	 	 else if (in[16:0] >= 231 && in <= 234) out = 2105;
	 	 	 else if (in[16:0] >= 235 && in <= 238) out = 2106;
	 	 	 else if (in[16:0] >= 239 && in <= 242) out = 2107;
	 	 	 else if (in[16:0] >= 243 && in <= 246) out = 2108;
	 	 	 else if (in[16:0] >= 247 && in <= 250) out = 2109;
	 	 	 else if (in[16:0] >= 251 && in <= 254) out = 2110;
	 	 	 else if (in[16:0] >= 255 && in <= 258) out = 2111;
	 	 	 else if (in[16:0] >= 259 && in <= 262) out = 2112;
	 	 	 else if (in[16:0] >= 263 && in <= 266) out = 2113;
	 	 	 else if (in[16:0] >= 267 && in <= 270) out = 2114;
	 	 	 else if (in[16:0] >= 271 && in <= 274) out = 2115;
	 	 	 else if (in[16:0] >= 275 && in <= 278) out = 2116;
	 	 	 else if (in[16:0] >= 279 && in <= 282) out = 2117;
	 	 	 else if (in[16:0] >= 283 && in <= 286) out = 2118;
	 	 	 else if (in[16:0] >= 287 && in <= 290) out = 2119;
	 	 	 else if (in[16:0] >= 291 && in <= 294) out = 2120;
	 	 	 else if (in[16:0] >= 295 && in <= 298) out = 2121;
	 	 	 else if (in[16:0] >= 299 && in <= 302) out = 2122;
	 	 	 else if (in[16:0] >= 303 && in <= 306) out = 2123;
	 	 	 else if (in[16:0] >= 307 && in <= 310) out = 2124;
	 	 	 else if (in[16:0] >= 311 && in <= 314) out = 2125;
	 	 	 else if (in[16:0] >= 315 && in <= 318) out = 2126;
	 	 	 else if (in[16:0] >= 319 && in <= 322) out = 2127;
	 	 	 else if (in[16:0] >= 323 && in <= 326) out = 2128;
	 	 	 else if (in[16:0] >= 327 && in <= 330) out = 2129;
	 	 	 else if (in[16:0] >= 331 && in <= 334) out = 2130;
	 	 	 else if (in[16:0] >= 335 && in <= 338) out = 2131;
	 	 	 else if (in[16:0] >= 339 && in <= 342) out = 2132;
	 	 	 else if (in[16:0] >= 343 && in <= 346) out = 2133;
	 	 	 else if (in[16:0] >= 347 && in <= 350) out = 2134;
	 	 	 else if (in[16:0] >= 351 && in <= 354) out = 2135;
	 	 	 else if (in[16:0] >= 355 && in <= 358) out = 2136;
	 	 	 else if (in[16:0] >= 359 && in <= 362) out = 2137;
	 	 	 else if (in[16:0] >= 363 && in <= 366) out = 2138;
	 	 	 else if (in[16:0] >= 367 && in <= 370) out = 2139;
	 	 	 else if (in[16:0] >= 371 && in <= 374) out = 2140;
	 	 	 else if (in[16:0] >= 375 && in <= 378) out = 2141;
	 	 	 else if (in[16:0] >= 379 && in <= 382) out = 2142;
	 	 	 else if (in[16:0] >= 383 && in <= 386) out = 2143;
	 	 	 else if (in[16:0] >= 387 && in <= 390) out = 2144;
	 	 	 else if (in[16:0] >= 391 && in <= 394) out = 2145;
	 	 	 else if (in[16:0] >= 395 && in <= 398) out = 2146;
	 	 	 else if (in[16:0] >= 399 && in <= 402) out = 2147;
	 	 	 else if (in[16:0] >= 403 && in <= 406) out = 2148;
	 	 	 else if (in[16:0] >= 407 && in <= 410) out = 2149;
	 	 	 else if (in[16:0] >= 411 && in <= 414) out = 2150;
	 	 	 else if (in[16:0] >= 415 && in <= 418) out = 2151;
	 	 	 else if (in[16:0] >= 419 && in <= 422) out = 2152;
	 	 	 else if (in[16:0] >= 423 && in <= 426) out = 2153;
	 	 	 else if (in[16:0] >= 427 && in <= 430) out = 2154;
	 	 	 else if (in[16:0] >= 431 && in <= 434) out = 2155;
	 	 	 else if (in[16:0] >= 435 && in <= 438) out = 2156;
	 	 	 else if (in[16:0] >= 439 && in <= 442) out = 2157;
	 	 	 else if (in[16:0] >= 443 && in <= 446) out = 2158;
	 	 	 else if (in[16:0] >= 447 && in <= 450) out = 2159;
	 	 	 else if (in[16:0] >= 451 && in <= 454) out = 2160;
	 	 	 else if (in[16:0] >= 455 && in <= 458) out = 2161;
	 	 	 else if (in[16:0] >= 459 && in <= 462) out = 2162;
	 	 	 else if (in[16:0] >= 463 && in <= 466) out = 2163;
	 	 	 else if (in[16:0] >= 467 && in <= 470) out = 2164;
	 	 	 else if (in[16:0] >= 471 && in <= 474) out = 2165;
	 	 	 else if (in[16:0] >= 475 && in <= 478) out = 2166;
	 	 	 else if (in[16:0] >= 479 && in <= 482) out = 2167;
	 	 	 else if (in[16:0] >= 483 && in <= 486) out = 2168;
	 	 	 else if (in[16:0] >= 487 && in <= 490) out = 2169;
	 	 	 else if (in[16:0] >= 491 && in <= 494) out = 2170;
	 	 	 else if (in[16:0] >= 495 && in <= 498) out = 2171;
	 	 	 else if (in[16:0] >= 499 && in <= 502) out = 2172;
	 	 	 else if (in[16:0] >= 503 && in <= 506) out = 2173;
	 	 	 else if (in[16:0] >= 507 && in <= 510) out = 2174;
	 	 	 else if (in[16:0] >= 511 && in <= 514) out = 2175;
	 	 	 else if (in[16:0] >= 515 && in <= 518) out = 2176;
	 	 	 else if (in[16:0] >= 519 && in <= 522) out = 2177;
	 	 	 else if (in[16:0] >= 523 && in <= 526) out = 2178;
	 	 	 else if (in[16:0] >= 527 && in <= 530) out = 2179;
	 	 	 else if (in[16:0] >= 531 && in <= 534) out = 2180;
	 	 	 else if (in[16:0] >= 535 && in <= 538) out = 2181;
	 	 	 else if (in[16:0] >= 539 && in <= 542) out = 2182;
	 	 	 else if (in[16:0] >= 543 && in <= 546) out = 2183;
	 	 	 else if (in[16:0] >= 547 && in <= 550) out = 2184;
	 	 	 else if (in[16:0] >= 551 && in <= 554) out = 2185;
	 	 	 else if (in[16:0] >= 555 && in <= 559) out = 2186;
	 	 	 else if (in[16:0] >= 560 && in <= 563) out = 2187;
	 	 	 else if (in[16:0] >= 564 && in <= 567) out = 2188;
	 	 	 else if (in[16:0] >= 568 && in <= 571) out = 2189;
	 	 	 else if (in[16:0] >= 572 && in <= 575) out = 2190;
	 	 	 else if (in[16:0] >= 576 && in <= 579) out = 2191;
	 	 	 else if (in[16:0] >= 580 && in <= 583) out = 2192;
	 	 	 else if (in[16:0] >= 584 && in <= 587) out = 2193;
	 	 	 else if (in[16:0] >= 588 && in <= 591) out = 2194;
	 	 	 else if (in[16:0] >= 592 && in <= 595) out = 2195;
	 	 	 else if (in[16:0] >= 596 && in <= 599) out = 2196;
	 	 	 else if (in[16:0] >= 600 && in <= 603) out = 2197;
	 	 	 else if (in[16:0] >= 604 && in <= 607) out = 2198;
	 	 	 else if (in[16:0] >= 608 && in <= 611) out = 2199;
	 	 	 else if (in[16:0] >= 612 && in <= 615) out = 2200;
	 	 	 else if (in[16:0] >= 616 && in <= 619) out = 2201;
	 	 	 else if (in[16:0] >= 620 && in <= 623) out = 2202;
	 	 	 else if (in[16:0] >= 624 && in <= 627) out = 2203;
	 	 	 else if (in[16:0] >= 628 && in <= 631) out = 2204;
	 	 	 else if (in[16:0] >= 632 && in <= 635) out = 2205;
	 	 	 else if (in[16:0] >= 636 && in <= 639) out = 2206;
	 	 	 else if (in[16:0] >= 640 && in <= 643) out = 2207;
	 	 	 else if (in[16:0] >= 644 && in <= 647) out = 2208;
	 	 	 else if (in[16:0] >= 648 && in <= 651) out = 2209;
	 	 	 else if (in[16:0] >= 652 && in <= 655) out = 2210;
	 	 	 else if (in[16:0] >= 656 && in <= 659) out = 2211;
	 	 	 else if (in[16:0] >= 660 && in <= 663) out = 2212;
	 	 	 else if (in[16:0] >= 664 && in <= 667) out = 2213;
	 	 	 else if (in[16:0] >= 668 && in <= 671) out = 2214;
	 	 	 else if (in[16:0] >= 672 && in <= 675) out = 2215;
	 	 	 else if (in[16:0] >= 676 && in <= 679) out = 2216;
	 	 	 else if (in[16:0] >= 680 && in <= 683) out = 2217;
	 	 	 else if (in[16:0] >= 684 && in <= 687) out = 2218;
	 	 	 else if (in[16:0] >= 688 && in <= 691) out = 2219;
	 	 	 else if (in[16:0] >= 692 && in <= 695) out = 2220;
	 	 	 else if (in[16:0] >= 696 && in <= 699) out = 2221;
	 	 	 else if (in[16:0] >= 700 && in <= 703) out = 2222;
	 	 	 else if (in[16:0] >= 704 && in <= 707) out = 2223;
	 	 	 else if (in[16:0] >= 708 && in <= 711) out = 2224;
	 	 	 else if (in[16:0] >= 712 && in <= 715) out = 2225;
	 	 	 else if (in[16:0] >= 716 && in <= 720) out = 2226;
	 	 	 else if (in[16:0] >= 721 && in <= 724) out = 2227;
	 	 	 else if (in[16:0] >= 725 && in <= 728) out = 2228;
	 	 	 else if (in[16:0] >= 729 && in <= 732) out = 2229;
	 	 	 else if (in[16:0] >= 733 && in <= 736) out = 2230;
	 	 	 else if (in[16:0] >= 737 && in <= 740) out = 2231;
	 	 	 else if (in[16:0] >= 741 && in <= 744) out = 2232;
	 	 	 else if (in[16:0] >= 745 && in <= 748) out = 2233;
	 	 	 else if (in[16:0] >= 749 && in <= 752) out = 2234;
	 	 	 else if (in[16:0] >= 753 && in <= 756) out = 2235;
	 	 	 else if (in[16:0] >= 757 && in <= 760) out = 2236;
	 	 	 else if (in[16:0] >= 761 && in <= 764) out = 2237;
	 	 	 else if (in[16:0] >= 765 && in <= 768) out = 2238;
	 	 	 else if (in[16:0] >= 769 && in <= 772) out = 2239;
	 	 	 else if (in[16:0] >= 773 && in <= 776) out = 2240;
	 	 	 else if (in[16:0] >= 777 && in <= 780) out = 2241;
	 	 	 else if (in[16:0] >= 781 && in <= 784) out = 2242;
	 	 	 else if (in[16:0] >= 785 && in <= 788) out = 2243;
	 	 	 else if (in[16:0] >= 789 && in <= 792) out = 2244;
	 	 	 else if (in[16:0] >= 793 && in <= 796) out = 2245;
	 	 	 else if (in[16:0] >= 797 && in <= 800) out = 2246;
	 	 	 else if (in[16:0] >= 801 && in <= 804) out = 2247;
	 	 	 else if (in[16:0] >= 805 && in <= 808) out = 2248;
	 	 	 else if (in[16:0] >= 809 && in <= 812) out = 2249;
	 	 	 else if (in[16:0] >= 813 && in <= 816) out = 2250;
	 	 	 else if (in[16:0] >= 817 && in <= 820) out = 2251;
	 	 	 else if (in[16:0] >= 821 && in <= 824) out = 2252;
	 	 	 else if (in[16:0] >= 825 && in <= 829) out = 2253;
	 	 	 else if (in[16:0] >= 830 && in <= 833) out = 2254;
	 	 	 else if (in[16:0] >= 834 && in <= 837) out = 2255;
	 	 	 else if (in[16:0] >= 838 && in <= 841) out = 2256;
	 	 	 else if (in[16:0] >= 842 && in <= 845) out = 2257;
	 	 	 else if (in[16:0] >= 846 && in <= 849) out = 2258;
	 	 	 else if (in[16:0] >= 850 && in <= 853) out = 2259;
	 	 	 else if (in[16:0] >= 854 && in <= 857) out = 2260;
	 	 	 else if (in[16:0] >= 858 && in <= 861) out = 2261;
	 	 	 else if (in[16:0] >= 862 && in <= 865) out = 2262;
	 	 	 else if (in[16:0] >= 866 && in <= 869) out = 2263;
	 	 	 else if (in[16:0] >= 870 && in <= 873) out = 2264;
	 	 	 else if (in[16:0] >= 874 && in <= 877) out = 2265;
	 	 	 else if (in[16:0] >= 878 && in <= 881) out = 2266;
	 	 	 else if (in[16:0] >= 882 && in <= 885) out = 2267;
	 	 	 else if (in[16:0] >= 886 && in <= 889) out = 2268;
	 	 	 else if (in[16:0] >= 890 && in <= 893) out = 2269;
	 	 	 else if (in[16:0] >= 894 && in <= 897) out = 2270;
	 	 	 else if (in[16:0] >= 898 && in <= 901) out = 2271;
	 	 	 else if (in[16:0] >= 902 && in <= 905) out = 2272;
	 	 	 else if (in[16:0] >= 906 && in <= 909) out = 2273;
	 	 	 else if (in[16:0] >= 910 && in <= 913) out = 2274;
	 	 	 else if (in[16:0] >= 914 && in <= 918) out = 2275;
	 	 	 else if (in[16:0] >= 919 && in <= 922) out = 2276;
	 	 	 else if (in[16:0] >= 923 && in <= 926) out = 2277;
	 	 	 else if (in[16:0] >= 927 && in <= 930) out = 2278;
	 	 	 else if (in[16:0] >= 931 && in <= 934) out = 2279;
	 	 	 else if (in[16:0] >= 935 && in <= 938) out = 2280;
	 	 	 else if (in[16:0] >= 939 && in <= 942) out = 2281;
	 	 	 else if (in[16:0] >= 943 && in <= 946) out = 2282;
	 	 	 else if (in[16:0] >= 947 && in <= 950) out = 2283;
	 	 	 else if (in[16:0] >= 951 && in <= 954) out = 2284;
	 	 	 else if (in[16:0] >= 955 && in <= 958) out = 2285;
	 	 	 else if (in[16:0] >= 959 && in <= 962) out = 2286;
	 	 	 else if (in[16:0] >= 963 && in <= 966) out = 2287;
	 	 	 else if (in[16:0] >= 967 && in <= 970) out = 2288;
	 	 	 else if (in[16:0] >= 971 && in <= 974) out = 2289;
	 	 	 else if (in[16:0] >= 975 && in <= 978) out = 2290;
	 	 	 else if (in[16:0] >= 979 && in <= 982) out = 2291;
	 	 	 else if (in[16:0] >= 983 && in <= 986) out = 2292;
	 	 	 else if (in[16:0] >= 987 && in <= 991) out = 2293;
	 	 	 else if (in[16:0] >= 992 && in <= 995) out = 2294;
	 	 	 else if (in[16:0] >= 996 && in <= 999) out = 2295;
	 	 	 else if (in[16:0] >= 1000 && in <= 1003) out = 2296;
	 	 	 else if (in[16:0] >= 1004 && in <= 1007) out = 2297;
	 	 	 else if (in[16:0] >= 1008 && in <= 1011) out = 2298;
	 	 	 else if (in[16:0] >= 1012 && in <= 1015) out = 2299;
	 	 	 else if (in[16:0] >= 1016 && in <= 1019) out = 2300;
	 	 	 else if (in[16:0] >= 1020 && in <= 1023) out = 2301;
	 	 	 else if (in[16:0] >= 1024 && in <= 1027) out = 2302;
	 	 	 else if (in[16:0] >= 1028 && in <= 1031) out = 2303;
	 	 	 else if (in[16:0] >= 1032 && in <= 1035) out = 2304;
	 	 	 else if (in[16:0] >= 1036 && in <= 1039) out = 2305;
	 	 	 else if (in[16:0] >= 1040 && in <= 1043) out = 2306;
	 	 	 else if (in[16:0] >= 1044 && in <= 1047) out = 2307;
	 	 	 else if (in[16:0] >= 1048 && in <= 1052) out = 2308;
	 	 	 else if (in[16:0] >= 1053 && in <= 1056) out = 2309;
	 	 	 else if (in[16:0] >= 1057 && in <= 1060) out = 2310;
	 	 	 else if (in[16:0] >= 1061 && in <= 1064) out = 2311;
	 	 	 else if (in[16:0] >= 1065 && in <= 1068) out = 2312;
	 	 	 else if (in[16:0] >= 1069 && in <= 1072) out = 2313;
	 	 	 else if (in[16:0] >= 1073 && in <= 1076) out = 2314;
	 	 	 else if (in[16:0] >= 1077 && in <= 1080) out = 2315;
	 	 	 else if (in[16:0] >= 1081 && in <= 1084) out = 2316;
	 	 	 else if (in[16:0] >= 1085 && in <= 1088) out = 2317;
	 	 	 else if (in[16:0] >= 1089 && in <= 1092) out = 2318;
	 	 	 else if (in[16:0] >= 1093 && in <= 1096) out = 2319;
	 	 	 else if (in[16:0] >= 1097 && in <= 1100) out = 2320;
	 	 	 else if (in[16:0] >= 1101 && in <= 1104) out = 2321;
	 	 	 else if (in[16:0] >= 1105 && in <= 1108) out = 2322;
	 	 	 else if (in[16:0] >= 1109 && in <= 1113) out = 2323;
	 	 	 else if (in[16:0] >= 1114 && in <= 1117) out = 2324;
	 	 	 else if (in[16:0] >= 1118 && in <= 1121) out = 2325;
	 	 	 else if (in[16:0] >= 1122 && in <= 1125) out = 2326;
	 	 	 else if (in[16:0] >= 1126 && in <= 1129) out = 2327;
	 	 	 else if (in[16:0] >= 1130 && in <= 1133) out = 2328;
	 	 	 else if (in[16:0] >= 1134 && in <= 1137) out = 2329;
	 	 	 else if (in[16:0] >= 1138 && in <= 1141) out = 2330;
	 	 	 else if (in[16:0] >= 1142 && in <= 1145) out = 2331;
	 	 	 else if (in[16:0] >= 1146 && in <= 1149) out = 2332;
	 	 	 else if (in[16:0] >= 1150 && in <= 1153) out = 2333;
	 	 	 else if (in[16:0] >= 1154 && in <= 1157) out = 2334;
	 	 	 else if (in[16:0] >= 1158 && in <= 1162) out = 2335;
	 	 	 else if (in[16:0] >= 1163 && in <= 1166) out = 2336;
	 	 	 else if (in[16:0] >= 1167 && in <= 1170) out = 2337;
	 	 	 else if (in[16:0] >= 1171 && in <= 1174) out = 2338;
	 	 	 else if (in[16:0] >= 1175 && in <= 1178) out = 2339;
	 	 	 else if (in[16:0] >= 1179 && in <= 1182) out = 2340;
	 	 	 else if (in[16:0] >= 1183 && in <= 1186) out = 2341;
	 	 	 else if (in[16:0] >= 1187 && in <= 1190) out = 2342;
	 	 	 else if (in[16:0] >= 1191 && in <= 1194) out = 2343;
	 	 	 else if (in[16:0] >= 1195 && in <= 1198) out = 2344;
	 	 	 else if (in[16:0] >= 1199 && in <= 1202) out = 2345;
	 	 	 else if (in[16:0] >= 1203 && in <= 1206) out = 2346;
	 	 	 else if (in[16:0] >= 1207 && in <= 1211) out = 2347;
	 	 	 else if (in[16:0] >= 1212 && in <= 1215) out = 2348;
	 	 	 else if (in[16:0] >= 1216 && in <= 1219) out = 2349;
	 	 	 else if (in[16:0] >= 1220 && in <= 1223) out = 2350;
	 	 	 else if (in[16:0] >= 1224 && in <= 1227) out = 2351;
	 	 	 else if (in[16:0] >= 1228 && in <= 1231) out = 2352;
	 	 	 else if (in[16:0] >= 1232 && in <= 1235) out = 2353;
	 	 	 else if (in[16:0] >= 1236 && in <= 1239) out = 2354;
	 	 	 else if (in[16:0] >= 1240 && in <= 1243) out = 2355;
	 	 	 else if (in[16:0] >= 1244 && in <= 1247) out = 2356;
	 	 	 else if (in[16:0] >= 1248 && in <= 1251) out = 2357;
	 	 	 else if (in[16:0] >= 1252 && in <= 1256) out = 2358;
	 	 	 else if (in[16:0] >= 1257 && in <= 1260) out = 2359;
	 	 	 else if (in[16:0] >= 1261 && in <= 1264) out = 2360;
	 	 	 else if (in[16:0] >= 1265 && in <= 1268) out = 2361;
	 	 	 else if (in[16:0] >= 1269 && in <= 1272) out = 2362;
	 	 	 else if (in[16:0] >= 1273 && in <= 1276) out = 2363;
	 	 	 else if (in[16:0] >= 1277 && in <= 1280) out = 2364;
	 	 	 else if (in[16:0] >= 1281 && in <= 1284) out = 2365;
	 	 	 else if (in[16:0] >= 1285 && in <= 1288) out = 2366;
	 	 	 else if (in[16:0] >= 1289 && in <= 1292) out = 2367;
	 	 	 else if (in[16:0] >= 1293 && in <= 1297) out = 2368;
	 	 	 else if (in[16:0] >= 1298 && in <= 1301) out = 2369;
	 	 	 else if (in[16:0] >= 1302 && in <= 1305) out = 2370;
	 	 	 else if (in[16:0] >= 1306 && in <= 1309) out = 2371;
	 	 	 else if (in[16:0] >= 1310 && in <= 1313) out = 2372;
	 	 	 else if (in[16:0] >= 1314 && in <= 1317) out = 2373;
	 	 	 else if (in[16:0] >= 1318 && in <= 1321) out = 2374;
	 	 	 else if (in[16:0] >= 1322 && in <= 1325) out = 2375;
	 	 	 else if (in[16:0] >= 1326 && in <= 1329) out = 2376;
	 	 	 else if (in[16:0] >= 1330 && in <= 1333) out = 2377;
	 	 	 else if (in[16:0] >= 1334 && in <= 1338) out = 2378;
	 	 	 else if (in[16:0] >= 1339 && in <= 1342) out = 2379;
	 	 	 else if (in[16:0] >= 1343 && in <= 1346) out = 2380;
	 	 	 else if (in[16:0] >= 1347 && in <= 1350) out = 2381;
	 	 	 else if (in[16:0] >= 1351 && in <= 1354) out = 2382;
	 	 	 else if (in[16:0] >= 1355 && in <= 1358) out = 2383;
	 	 	 else if (in[16:0] >= 1359 && in <= 1362) out = 2384;
	 	 	 else if (in[16:0] >= 1363 && in <= 1366) out = 2385;
	 	 	 else if (in[16:0] >= 1367 && in <= 1370) out = 2386;
	 	 	 else if (in[16:0] >= 1371 && in <= 1375) out = 2387;
	 	 	 else if (in[16:0] >= 1376 && in <= 1379) out = 2388;
	 	 	 else if (in[16:0] >= 1380 && in <= 1383) out = 2389;
	 	 	 else if (in[16:0] >= 1384 && in <= 1387) out = 2390;
	 	 	 else if (in[16:0] >= 1388 && in <= 1391) out = 2391;
	 	 	 else if (in[16:0] >= 1392 && in <= 1395) out = 2392;
	 	 	 else if (in[16:0] >= 1396 && in <= 1399) out = 2393;
	 	 	 else if (in[16:0] >= 1400 && in <= 1403) out = 2394;
	 	 	 else if (in[16:0] >= 1404 && in <= 1408) out = 2395;
	 	 	 else if (in[16:0] >= 1409 && in <= 1412) out = 2396;
	 	 	 else if (in[16:0] >= 1413 && in <= 1416) out = 2397;
	 	 	 else if (in[16:0] >= 1417 && in <= 1420) out = 2398;
	 	 	 else if (in[16:0] >= 1421 && in <= 1424) out = 2399;
	 	 	 else if (in[16:0] >= 1425 && in <= 1428) out = 2400;
	 	 	 else if (in[16:0] >= 1429 && in <= 1432) out = 2401;
	 	 	 else if (in[16:0] >= 1433 && in <= 1436) out = 2402;
	 	 	 else if (in[16:0] >= 1437 && in <= 1441) out = 2403;
	 	 	 else if (in[16:0] >= 1442 && in <= 1445) out = 2404;
	 	 	 else if (in[16:0] >= 1446 && in <= 1449) out = 2405;
	 	 	 else if (in[16:0] >= 1450 && in <= 1453) out = 2406;
	 	 	 else if (in[16:0] >= 1454 && in <= 1457) out = 2407;
	 	 	 else if (in[16:0] >= 1458 && in <= 1461) out = 2408;
	 	 	 else if (in[16:0] >= 1462 && in <= 1465) out = 2409;
	 	 	 else if (in[16:0] >= 1466 && in <= 1469) out = 2410;
	 	 	 else if (in[16:0] >= 1470 && in <= 1474) out = 2411;
	 	 	 else if (in[16:0] >= 1475 && in <= 1478) out = 2412;
	 	 	 else if (in[16:0] >= 1479 && in <= 1482) out = 2413;
	 	 	 else if (in[16:0] >= 1483 && in <= 1486) out = 2414;
	 	 	 else if (in[16:0] >= 1487 && in <= 1490) out = 2415;
	 	 	 else if (in[16:0] >= 1491 && in <= 1494) out = 2416;
	 	 	 else if (in[16:0] >= 1495 && in <= 1498) out = 2417;
	 	 	 else if (in[16:0] >= 1499 && in <= 1503) out = 2418;
	 	 	 else if (in[16:0] >= 1504 && in <= 1507) out = 2419;
	 	 	 else if (in[16:0] >= 1508 && in <= 1511) out = 2420;
	 	 	 else if (in[16:0] >= 1512 && in <= 1515) out = 2421;
	 	 	 else if (in[16:0] >= 1516 && in <= 1519) out = 2422;
	 	 	 else if (in[16:0] >= 1520 && in <= 1523) out = 2423;
	 	 	 else if (in[16:0] >= 1524 && in <= 1527) out = 2424;
	 	 	 else if (in[16:0] >= 1528 && in <= 1531) out = 2425;
	 	 	 else if (in[16:0] >= 1532 && in <= 1536) out = 2426;
	 	 	 else if (in[16:0] >= 1537 && in <= 1540) out = 2427;
	 	 	 else if (in[16:0] >= 1541 && in <= 1544) out = 2428;
	 	 	 else if (in[16:0] >= 1545 && in <= 1548) out = 2429;
	 	 	 else if (in[16:0] >= 1549 && in <= 1552) out = 2430;
	 	 	 else if (in[16:0] >= 1553 && in <= 1556) out = 2431;
	 	 	 else if (in[16:0] >= 1557 && in <= 1560) out = 2432;
	 	 	 else if (in[16:0] >= 1561 && in <= 1565) out = 2433;
	 	 	 else if (in[16:0] >= 1566 && in <= 1569) out = 2434;
	 	 	 else if (in[16:0] >= 1570 && in <= 1573) out = 2435;
	 	 	 else if (in[16:0] >= 1574 && in <= 1577) out = 2436;
	 	 	 else if (in[16:0] >= 1578 && in <= 1581) out = 2437;
	 	 	 else if (in[16:0] >= 1582 && in <= 1585) out = 2438;
	 	 	 else if (in[16:0] >= 1586 && in <= 1590) out = 2439;
	 	 	 else if (in[16:0] >= 1591 && in <= 1594) out = 2440;
	 	 	 else if (in[16:0] >= 1595 && in <= 1598) out = 2441;
	 	 	 else if (in[16:0] >= 1599 && in <= 1602) out = 2442;
	 	 	 else if (in[16:0] >= 1603 && in <= 1606) out = 2443;
	 	 	 else if (in[16:0] >= 1607 && in <= 1610) out = 2444;
	 	 	 else if (in[16:0] >= 1611 && in <= 1614) out = 2445;
	 	 	 else if (in[16:0] >= 1615 && in <= 1619) out = 2446;
	 	 	 else if (in[16:0] >= 1620 && in <= 1623) out = 2447;
	 	 	 else if (in[16:0] >= 1624 && in <= 1627) out = 2448;
	 	 	 else if (in[16:0] >= 1628 && in <= 1631) out = 2449;
	 	 	 else if (in[16:0] >= 1632 && in <= 1635) out = 2450;
	 	 	 else if (in[16:0] >= 1636 && in <= 1639) out = 2451;
	 	 	 else if (in[16:0] >= 1640 && in <= 1644) out = 2452;
	 	 	 else if (in[16:0] >= 1645 && in <= 1648) out = 2453;
	 	 	 else if (in[16:0] >= 1649 && in <= 1652) out = 2454;
	 	 	 else if (in[16:0] >= 1653 && in <= 1656) out = 2455;
	 	 	 else if (in[16:0] >= 1657 && in <= 1660) out = 2456;
	 	 	 else if (in[16:0] >= 1661 && in <= 1664) out = 2457;
	 	 	 else if (in[16:0] >= 1665 && in <= 1669) out = 2458;
	 	 	 else if (in[16:0] >= 1670 && in <= 1673) out = 2459;
	 	 	 else if (in[16:0] >= 1674 && in <= 1677) out = 2460;
	 	 	 else if (in[16:0] >= 1678 && in <= 1681) out = 2461;
	 	 	 else if (in[16:0] >= 1682 && in <= 1685) out = 2462;
	 	 	 else if (in[16:0] >= 1686 && in <= 1689) out = 2463;
	 	 	 else if (in[16:0] >= 1690 && in <= 1694) out = 2464;
	 	 	 else if (in[16:0] >= 1695 && in <= 1698) out = 2465;
	 	 	 else if (in[16:0] >= 1699 && in <= 1702) out = 2466;
	 	 	 else if (in[16:0] >= 1703 && in <= 1706) out = 2467;
	 	 	 else if (in[16:0] >= 1707 && in <= 1710) out = 2468;
	 	 	 else if (in[16:0] >= 1711 && in <= 1715) out = 2469;
	 	 	 else if (in[16:0] >= 1716 && in <= 1719) out = 2470;
	 	 	 else if (in[16:0] >= 1720 && in <= 1723) out = 2471;
	 	 	 else if (in[16:0] >= 1724 && in <= 1727) out = 2472;
	 	 	 else if (in[16:0] >= 1728 && in <= 1731) out = 2473;
	 	 	 else if (in[16:0] >= 1732 && in <= 1735) out = 2474;
	 	 	 else if (in[16:0] >= 1736 && in <= 1740) out = 2475;
	 	 	 else if (in[16:0] >= 1741 && in <= 1744) out = 2476;
	 	 	 else if (in[16:0] >= 1745 && in <= 1748) out = 2477;
	 	 	 else if (in[16:0] >= 1749 && in <= 1752) out = 2478;
	 	 	 else if (in[16:0] >= 1753 && in <= 1756) out = 2479;
	 	 	 else if (in[16:0] >= 1757 && in <= 1761) out = 2480;
	 	 	 else if (in[16:0] >= 1762 && in <= 1765) out = 2481;
	 	 	 else if (in[16:0] >= 1766 && in <= 1769) out = 2482;
	 	 	 else if (in[16:0] >= 1770 && in <= 1773) out = 2483;
	 	 	 else if (in[16:0] >= 1774 && in <= 1777) out = 2484;
	 	 	 else if (in[16:0] >= 1778 && in <= 1782) out = 2485;
	 	 	 else if (in[16:0] >= 1783 && in <= 1786) out = 2486;
	 	 	 else if (in[16:0] >= 1787 && in <= 1790) out = 2487;
	 	 	 else if (in[16:0] >= 1791 && in <= 1794) out = 2488;
	 	 	 else if (in[16:0] >= 1795 && in <= 1798) out = 2489;
	 	 	 else if (in[16:0] >= 1799 && in <= 1802) out = 2490;
	 	 	 else if (in[16:0] >= 1803 && in <= 1807) out = 2491;
	 	 	 else if (in[16:0] >= 1808 && in <= 1811) out = 2492;
	 	 	 else if (in[16:0] >= 1812 && in <= 1815) out = 2493;
	 	 	 else if (in[16:0] >= 1816 && in <= 1819) out = 2494;
	 	 	 else if (in[16:0] >= 1820 && in <= 1823) out = 2495;
	 	 	 else if (in[16:0] >= 1824 && in <= 1828) out = 2496;
	 	 	 else if (in[16:0] >= 1829 && in <= 1832) out = 2497;
	 	 	 else if (in[16:0] >= 1833 && in <= 1836) out = 2498;
	 	 	 else if (in[16:0] >= 1837 && in <= 1840) out = 2499;
	 	 	 else if (in[16:0] >= 1841 && in <= 1845) out = 2500;
	 	 	 else if (in[16:0] >= 1846 && in <= 1849) out = 2501;
	 	 	 else if (in[16:0] >= 1850 && in <= 1853) out = 2502;
	 	 	 else if (in[16:0] >= 1854 && in <= 1857) out = 2503;
	 	 	 else if (in[16:0] >= 1858 && in <= 1861) out = 2504;
	 	 	 else if (in[16:0] >= 1862 && in <= 1866) out = 2505;
	 	 	 else if (in[16:0] >= 1867 && in <= 1870) out = 2506;
	 	 	 else if (in[16:0] >= 1871 && in <= 1874) out = 2507;
	 	 	 else if (in[16:0] >= 1875 && in <= 1878) out = 2508;
	 	 	 else if (in[16:0] >= 1879 && in <= 1882) out = 2509;
	 	 	 else if (in[16:0] >= 1883 && in <= 1887) out = 2510;
	 	 	 else if (in[16:0] >= 1888 && in <= 1891) out = 2511;
	 	 	 else if (in[16:0] >= 1892 && in <= 1895) out = 2512;
	 	 	 else if (in[16:0] >= 1896 && in <= 1899) out = 2513;
	 	 	 else if (in[16:0] >= 1900 && in <= 1904) out = 2514;
	 	 	 else if (in[16:0] >= 1905 && in <= 1908) out = 2515;
	 	 	 else if (in[16:0] >= 1909 && in <= 1912) out = 2516;
	 	 	 else if (in[16:0] >= 1913 && in <= 1916) out = 2517;
	 	 	 else if (in[16:0] >= 1917 && in <= 1920) out = 2518;
	 	 	 else if (in[16:0] >= 1921 && in <= 1925) out = 2519;
	 	 	 else if (in[16:0] >= 1926 && in <= 1929) out = 2520;
	 	 	 else if (in[16:0] >= 1930 && in <= 1933) out = 2521;
	 	 	 else if (in[16:0] >= 1934 && in <= 1937) out = 2522;
	 	 	 else if (in[16:0] >= 1938 && in <= 1942) out = 2523;
	 	 	 else if (in[16:0] >= 1943 && in <= 1946) out = 2524;
	 	 	 else if (in[16:0] >= 1947 && in <= 1950) out = 2525;
	 	 	 else if (in[16:0] >= 1951 && in <= 1954) out = 2526;
	 	 	 else if (in[16:0] >= 1955 && in <= 1958) out = 2527;
	 	 	 else if (in[16:0] >= 1959 && in <= 1963) out = 2528;
	 	 	 else if (in[16:0] >= 1964 && in <= 1967) out = 2529;
	 	 	 else if (in[16:0] >= 1968 && in <= 1971) out = 2530;
	 	 	 else if (in[16:0] >= 1972 && in <= 1975) out = 2531;
	 	 	 else if (in[16:0] >= 1976 && in <= 1980) out = 2532;
	 	 	 else if (in[16:0] >= 1981 && in <= 1984) out = 2533;
	 	 	 else if (in[16:0] >= 1985 && in <= 1988) out = 2534;
	 	 	 else if (in[16:0] >= 1989 && in <= 1992) out = 2535;
	 	 	 else if (in[16:0] >= 1993 && in <= 1997) out = 2536;
	 	 	 else if (in[16:0] >= 1998 && in <= 2001) out = 2537;
	 	 	 else if (in[16:0] >= 2002 && in <= 2005) out = 2538;
	 	 	 else if (in[16:0] >= 2006 && in <= 2009) out = 2539;
	 	 	 else if (in[16:0] >= 2010 && in <= 2014) out = 2540;
	 	 	 else if (in[16:0] >= 2015 && in <= 2018) out = 2541;
	 	 	 else if (in[16:0] >= 2019 && in <= 2022) out = 2542;
	 	 	 else if (in[16:0] >= 2023 && in <= 2026) out = 2543;
	 	 	 else if (in[16:0] >= 2027 && in <= 2031) out = 2544;
	 	 	 else if (in[16:0] >= 2032 && in <= 2035) out = 2545;
	 	 	 else if (in[16:0] >= 2036 && in <= 2039) out = 2546;
	 	 	 else if (in[16:0] >= 2040 && in <= 2043) out = 2547;
	 	 	 else if (in[16:0] >= 2044 && in <= 2048) out = 2548;
	 	 	 else if (in[16:0] >= 2049 && in <= 2052) out = 2549;
	 	 	 else if (in[16:0] >= 2053 && in <= 2056) out = 2550;
	 	 	 else if (in[16:0] >= 2057 && in <= 2060) out = 2551;
	 	 	 else if (in[16:0] >= 2061 && in <= 2065) out = 2552;
	 	 	 else if (in[16:0] >= 2066 && in <= 2069) out = 2553;
	 	 	 else if (in[16:0] >= 2070 && in <= 2073) out = 2554;
	 	 	 else if (in[16:0] >= 2074 && in <= 2077) out = 2555;
	 	 	 else if (in[16:0] >= 2078 && in <= 2082) out = 2556;
	 	 	 else if (in[16:0] >= 2083 && in <= 2086) out = 2557;
	 	 	 else if (in[16:0] >= 2087 && in <= 2090) out = 2558;
	 	 	 else if (in[16:0] >= 2091 && in <= 2095) out = 2559;
	 	 	 else if (in[16:0] >= 2096 && in <= 2099) out = 2560;
	 	 	 else if (in[16:0] >= 2100 && in <= 2103) out = 2561;
	 	 	 else if (in[16:0] >= 2104 && in <= 2107) out = 2562;
	 	 	 else if (in[16:0] >= 2108 && in <= 2112) out = 2563;
	 	 	 else if (in[16:0] >= 2113 && in <= 2116) out = 2564;
	 	 	 else if (in[16:0] >= 2117 && in <= 2120) out = 2565;
	 	 	 else if (in[16:0] >= 2121 && in <= 2124) out = 2566;
	 	 	 else if (in[16:0] >= 2125 && in <= 2129) out = 2567;
	 	 	 else if (in[16:0] >= 2130 && in <= 2133) out = 2568;
	 	 	 else if (in[16:0] >= 2134 && in <= 2137) out = 2569;
	 	 	 else if (in[16:0] >= 2138 && in <= 2142) out = 2570;
	 	 	 else if (in[16:0] >= 2143 && in <= 2146) out = 2571;
	 	 	 else if (in[16:0] >= 2147 && in <= 2150) out = 2572;
	 	 	 else if (in[16:0] >= 2151 && in <= 2154) out = 2573;
	 	 	 else if (in[16:0] >= 2155 && in <= 2159) out = 2574;
	 	 	 else if (in[16:0] >= 2160 && in <= 2163) out = 2575;
	 	 	 else if (in[16:0] >= 2164 && in <= 2167) out = 2576;
	 	 	 else if (in[16:0] >= 2168 && in <= 2172) out = 2577;
	 	 	 else if (in[16:0] >= 2173 && in <= 2176) out = 2578;
	 	 	 else if (in[16:0] >= 2177 && in <= 2180) out = 2579;
	 	 	 else if (in[16:0] >= 2181 && in <= 2184) out = 2580;
	 	 	 else if (in[16:0] >= 2185 && in <= 2189) out = 2581;
	 	 	 else if (in[16:0] >= 2190 && in <= 2193) out = 2582;
	 	 	 else if (in[16:0] >= 2194 && in <= 2197) out = 2583;
	 	 	 else if (in[16:0] >= 2198 && in <= 2202) out = 2584;
	 	 	 else if (in[16:0] >= 2203 && in <= 2206) out = 2585;
	 	 	 else if (in[16:0] >= 2207 && in <= 2210) out = 2586;
	 	 	 else if (in[16:0] >= 2211 && in <= 2214) out = 2587;
	 	 	 else if (in[16:0] >= 2215 && in <= 2219) out = 2588;
	 	 	 else if (in[16:0] >= 2220 && in <= 2223) out = 2589;
	 	 	 else if (in[16:0] >= 2224 && in <= 2227) out = 2590;
	 	 	 else if (in[16:0] >= 2228 && in <= 2232) out = 2591;
	 	 	 else if (in[16:0] >= 2233 && in <= 2236) out = 2592;
	 	 	 else if (in[16:0] >= 2237 && in <= 2240) out = 2593;
	 	 	 else if (in[16:0] >= 2241 && in <= 2245) out = 2594;
	 	 	 else if (in[16:0] >= 2246 && in <= 2249) out = 2595;
	 	 	 else if (in[16:0] >= 2250 && in <= 2253) out = 2596;
	 	 	 else if (in[16:0] >= 2254 && in <= 2258) out = 2597;
	 	 	 else if (in[16:0] >= 2259 && in <= 2262) out = 2598;
	 	 	 else if (in[16:0] >= 2263 && in <= 2266) out = 2599;
	 	 	 else if (in[16:0] >= 2267 && in <= 2270) out = 2600;
	 	 	 else if (in[16:0] >= 2271 && in <= 2275) out = 2601;
	 	 	 else if (in[16:0] >= 2276 && in <= 2279) out = 2602;
	 	 	 else if (in[16:0] >= 2280 && in <= 2283) out = 2603;
	 	 	 else if (in[16:0] >= 2284 && in <= 2288) out = 2604;
	 	 	 else if (in[16:0] >= 2289 && in <= 2292) out = 2605;
	 	 	 else if (in[16:0] >= 2293 && in <= 2296) out = 2606;
	 	 	 else if (in[16:0] >= 2297 && in <= 2301) out = 2607;
	 	 	 else if (in[16:0] >= 2302 && in <= 2305) out = 2608;
	 	 	 else if (in[16:0] >= 2306 && in <= 2309) out = 2609;
	 	 	 else if (in[16:0] >= 2310 && in <= 2314) out = 2610;
	 	 	 else if (in[16:0] >= 2315 && in <= 2318) out = 2611;
	 	 	 else if (in[16:0] >= 2319 && in <= 2322) out = 2612;
	 	 	 else if (in[16:0] >= 2323 && in <= 2327) out = 2613;
	 	 	 else if (in[16:0] >= 2328 && in <= 2331) out = 2614;
	 	 	 else if (in[16:0] >= 2332 && in <= 2335) out = 2615;
	 	 	 else if (in[16:0] >= 2336 && in <= 2340) out = 2616;
	 	 	 else if (in[16:0] >= 2341 && in <= 2344) out = 2617;
	 	 	 else if (in[16:0] >= 2345 && in <= 2348) out = 2618;
	 	 	 else if (in[16:0] >= 2349 && in <= 2353) out = 2619;
	 	 	 else if (in[16:0] >= 2354 && in <= 2357) out = 2620;
	 	 	 else if (in[16:0] >= 2358 && in <= 2361) out = 2621;
	 	 	 else if (in[16:0] >= 2362 && in <= 2366) out = 2622;
	 	 	 else if (in[16:0] >= 2367 && in <= 2370) out = 2623;
	 	 	 else if (in[16:0] >= 2371 && in <= 2374) out = 2624;
	 	 	 else if (in[16:0] >= 2375 && in <= 2379) out = 2625;
	 	 	 else if (in[16:0] >= 2380 && in <= 2383) out = 2626;
	 	 	 else if (in[16:0] >= 2384 && in <= 2387) out = 2627;
	 	 	 else if (in[16:0] >= 2388 && in <= 2392) out = 2628;
	 	 	 else if (in[16:0] >= 2393 && in <= 2396) out = 2629;
	 	 	 else if (in[16:0] >= 2397 && in <= 2401) out = 2630;
	 	 	 else if (in[16:0] >= 2402 && in <= 2405) out = 2631;
	 	 	 else if (in[16:0] >= 2406 && in <= 2409) out = 2632;
	 	 	 else if (in[16:0] >= 2410 && in <= 2414) out = 2633;
	 	 	 else if (in[16:0] >= 2415 && in <= 2418) out = 2634;
	 	 	 else if (in[16:0] >= 2419 && in <= 2422) out = 2635;
	 	 	 else if (in[16:0] >= 2423 && in <= 2427) out = 2636;
	 	 	 else if (in[16:0] >= 2428 && in <= 2431) out = 2637;
	 	 	 else if (in[16:0] >= 2432 && in <= 2435) out = 2638;
	 	 	 else if (in[16:0] >= 2436 && in <= 2440) out = 2639;
	 	 	 else if (in[16:0] >= 2441 && in <= 2444) out = 2640;
	 	 	 else if (in[16:0] >= 2445 && in <= 2449) out = 2641;
	 	 	 else if (in[16:0] >= 2450 && in <= 2453) out = 2642;
	 	 	 else if (in[16:0] >= 2454 && in <= 2457) out = 2643;
	 	 	 else if (in[16:0] >= 2458 && in <= 2462) out = 2644;
	 	 	 else if (in[16:0] >= 2463 && in <= 2466) out = 2645;
	 	 	 else if (in[16:0] >= 2467 && in <= 2470) out = 2646;
	 	 	 else if (in[16:0] >= 2471 && in <= 2475) out = 2647;
	 	 	 else if (in[16:0] >= 2476 && in <= 2479) out = 2648;
	 	 	 else if (in[16:0] >= 2480 && in <= 2484) out = 2649;
	 	 	 else if (in[16:0] >= 2485 && in <= 2488) out = 2650;
	 	 	 else if (in[16:0] >= 2489 && in <= 2492) out = 2651;
	 	 	 else if (in[16:0] >= 2493 && in <= 2497) out = 2652;
	 	 	 else if (in[16:0] >= 2498 && in <= 2501) out = 2653;
	 	 	 else if (in[16:0] >= 2502 && in <= 2505) out = 2654;
	 	 	 else if (in[16:0] >= 2506 && in <= 2510) out = 2655;
	 	 	 else if (in[16:0] >= 2511 && in <= 2514) out = 2656;
	 	 	 else if (in[16:0] >= 2515 && in <= 2519) out = 2657;
	 	 	 else if (in[16:0] >= 2520 && in <= 2523) out = 2658;
	 	 	 else if (in[16:0] >= 2524 && in <= 2527) out = 2659;
	 	 	 else if (in[16:0] >= 2528 && in <= 2532) out = 2660;
	 	 	 else if (in[16:0] >= 2533 && in <= 2536) out = 2661;
	 	 	 else if (in[16:0] >= 2537 && in <= 2541) out = 2662;
	 	 	 else if (in[16:0] >= 2542 && in <= 2545) out = 2663;
	 	 	 else if (in[16:0] >= 2546 && in <= 2549) out = 2664;
	 	 	 else if (in[16:0] >= 2550 && in <= 2554) out = 2665;
	 	 	 else if (in[16:0] >= 2555 && in <= 2558) out = 2666;
	 	 	 else if (in[16:0] >= 2559 && in <= 2563) out = 2667;
	 	 	 else if (in[16:0] >= 2564 && in <= 2567) out = 2668;
	 	 	 else if (in[16:0] >= 2568 && in <= 2571) out = 2669;
	 	 	 else if (in[16:0] >= 2572 && in <= 2576) out = 2670;
	 	 	 else if (in[16:0] >= 2577 && in <= 2580) out = 2671;
	 	 	 else if (in[16:0] >= 2581 && in <= 2585) out = 2672;
	 	 	 else if (in[16:0] >= 2586 && in <= 2589) out = 2673;
	 	 	 else if (in[16:0] >= 2590 && in <= 2593) out = 2674;
	 	 	 else if (in[16:0] >= 2594 && in <= 2598) out = 2675;
	 	 	 else if (in[16:0] >= 2599 && in <= 2602) out = 2676;
	 	 	 else if (in[16:0] >= 2603 && in <= 2607) out = 2677;
	 	 	 else if (in[16:0] >= 2608 && in <= 2611) out = 2678;
	 	 	 else if (in[16:0] >= 2612 && in <= 2616) out = 2679;
	 	 	 else if (in[16:0] >= 2617 && in <= 2620) out = 2680;
	 	 	 else if (in[16:0] >= 2621 && in <= 2624) out = 2681;
	 	 	 else if (in[16:0] >= 2625 && in <= 2629) out = 2682;
	 	 	 else if (in[16:0] >= 2630 && in <= 2633) out = 2683;
	 	 	 else if (in[16:0] >= 2634 && in <= 2638) out = 2684;
	 	 	 else if (in[16:0] >= 2639 && in <= 2642) out = 2685;
	 	 	 else if (in[16:0] >= 2643 && in <= 2647) out = 2686;
	 	 	 else if (in[16:0] >= 2648 && in <= 2651) out = 2687;
	 	 	 else if (in[16:0] >= 2652 && in <= 2655) out = 2688;
	 	 	 else if (in[16:0] >= 2656 && in <= 2660) out = 2689;
	 	 	 else if (in[16:0] >= 2661 && in <= 2664) out = 2690;
	 	 	 else if (in[16:0] >= 2665 && in <= 2669) out = 2691;
	 	 	 else if (in[16:0] >= 2670 && in <= 2673) out = 2692;
	 	 	 else if (in[16:0] >= 2674 && in <= 2678) out = 2693;
	 	 	 else if (in[16:0] >= 2679 && in <= 2682) out = 2694;
	 	 	 else if (in[16:0] >= 2683 && in <= 2687) out = 2695;
	 	 	 else if (in[16:0] >= 2688 && in <= 2691) out = 2696;
	 	 	 else if (in[16:0] >= 2692 && in <= 2695) out = 2697;
	 	 	 else if (in[16:0] >= 2696 && in <= 2700) out = 2698;
	 	 	 else if (in[16:0] >= 2701 && in <= 2704) out = 2699;
	 	 	 else if (in[16:0] >= 2705 && in <= 2709) out = 2700;
	 	 	 else if (in[16:0] >= 2710 && in <= 2713) out = 2701;
	 	 	 else if (in[16:0] >= 2714 && in <= 2718) out = 2702;
	 	 	 else if (in[16:0] >= 2719 && in <= 2722) out = 2703;
	 	 	 else if (in[16:0] >= 2723 && in <= 2727) out = 2704;
	 	 	 else if (in[16:0] >= 2728 && in <= 2731) out = 2705;
	 	 	 else if (in[16:0] >= 2732 && in <= 2736) out = 2706;
	 	 	 else if (in[16:0] >= 2737 && in <= 2740) out = 2707;
	 	 	 else if (in[16:0] >= 2741 && in <= 2744) out = 2708;
	 	 	 else if (in[16:0] >= 2745 && in <= 2749) out = 2709;
	 	 	 else if (in[16:0] >= 2750 && in <= 2753) out = 2710;
	 	 	 else if (in[16:0] >= 2754 && in <= 2758) out = 2711;
	 	 	 else if (in[16:0] >= 2759 && in <= 2762) out = 2712;
	 	 	 else if (in[16:0] >= 2763 && in <= 2767) out = 2713;
	 	 	 else if (in[16:0] >= 2768 && in <= 2771) out = 2714;
	 	 	 else if (in[16:0] >= 2772 && in <= 2776) out = 2715;
	 	 	 else if (in[16:0] >= 2777 && in <= 2780) out = 2716;
	 	 	 else if (in[16:0] >= 2781 && in <= 2785) out = 2717;
	 	 	 else if (in[16:0] >= 2786 && in <= 2789) out = 2718;
	 	 	 else if (in[16:0] >= 2790 && in <= 2794) out = 2719;
	 	 	 else if (in[16:0] >= 2795 && in <= 2798) out = 2720;
	 	 	 else if (in[16:0] >= 2799 && in <= 2803) out = 2721;
	 	 	 else if (in[16:0] >= 2804 && in <= 2807) out = 2722;
	 	 	 else if (in[16:0] >= 2808 && in <= 2812) out = 2723;
	 	 	 else if (in[16:0] >= 2813 && in <= 2816) out = 2724;
	 	 	 else if (in[16:0] >= 2817 && in <= 2821) out = 2725;
	 	 	 else if (in[16:0] >= 2822 && in <= 2825) out = 2726;
	 	 	 else if (in[16:0] >= 2826 && in <= 2830) out = 2727;
	 	 	 else if (in[16:0] >= 2831 && in <= 2834) out = 2728;
	 	 	 else if (in[16:0] >= 2835 && in <= 2839) out = 2729;
	 	 	 else if (in[16:0] >= 2840 && in <= 2843) out = 2730;
	 	 	 else if (in[16:0] >= 2844 && in <= 2848) out = 2731;
	 	 	 else if (in[16:0] >= 2849 && in <= 2852) out = 2732;
	 	 	 else if (in[16:0] >= 2853 && in <= 2857) out = 2733;
	 	 	 else if (in[16:0] >= 2858 && in <= 2861) out = 2734;
	 	 	 else if (in[16:0] >= 2862 && in <= 2866) out = 2735;
	 	 	 else if (in[16:0] >= 2867 && in <= 2870) out = 2736;
	 	 	 else if (in[16:0] >= 2871 && in <= 2875) out = 2737;
	 	 	 else if (in[16:0] >= 2876 && in <= 2879) out = 2738;
	 	 	 else if (in[16:0] >= 2880 && in <= 2884) out = 2739;
	 	 	 else if (in[16:0] >= 2885 && in <= 2888) out = 2740;
	 	 	 else if (in[16:0] >= 2889 && in <= 2893) out = 2741;
	 	 	 else if (in[16:0] >= 2894 && in <= 2897) out = 2742;
	 	 	 else if (in[16:0] >= 2898 && in <= 2902) out = 2743;
	 	 	 else if (in[16:0] >= 2903 && in <= 2906) out = 2744;
	 	 	 else if (in[16:0] >= 2907 && in <= 2911) out = 2745;
	 	 	 else if (in[16:0] >= 2912 && in <= 2915) out = 2746;
	 	 	 else if (in[16:0] >= 2916 && in <= 2920) out = 2747;
	 	 	 else if (in[16:0] >= 2921 && in <= 2924) out = 2748;
	 	 	 else if (in[16:0] >= 2925 && in <= 2929) out = 2749;
	 	 	 else if (in[16:0] >= 2930 && in <= 2934) out = 2750;
	 	 	 else if (in[16:0] >= 2935 && in <= 2938) out = 2751;
	 	 	 else if (in[16:0] >= 2939 && in <= 2943) out = 2752;
	 	 	 else if (in[16:0] >= 2944 && in <= 2947) out = 2753;
	 	 	 else if (in[16:0] >= 2948 && in <= 2952) out = 2754;
	 	 	 else if (in[16:0] >= 2953 && in <= 2956) out = 2755;
	 	 	 else if (in[16:0] >= 2957 && in <= 2961) out = 2756;
	 	 	 else if (in[16:0] >= 2962 && in <= 2965) out = 2757;
	 	 	 else if (in[16:0] >= 2966 && in <= 2970) out = 2758;
	 	 	 else if (in[16:0] >= 2971 && in <= 2974) out = 2759;
	 	 	 else if (in[16:0] >= 2975 && in <= 2979) out = 2760;
	 	 	 else if (in[16:0] >= 2980 && in <= 2984) out = 2761;
	 	 	 else if (in[16:0] >= 2985 && in <= 2988) out = 2762;
	 	 	 else if (in[16:0] >= 2989 && in <= 2993) out = 2763;
	 	 	 else if (in[16:0] >= 2994 && in <= 2997) out = 2764;
	 	 	 else if (in[16:0] >= 2998 && in <= 3002) out = 2765;
	 	 	 else if (in[16:0] >= 3003 && in <= 3006) out = 2766;
	 	 	 else if (in[16:0] >= 3007 && in <= 3011) out = 2767;
	 	 	 else if (in[16:0] >= 3012 && in <= 3015) out = 2768;
	 	 	 else if (in[16:0] >= 3016 && in <= 3020) out = 2769;
	 	 	 else if (in[16:0] >= 3021 && in <= 3025) out = 2770;
	 	 	 else if (in[16:0] >= 3026 && in <= 3029) out = 2771;
	 	 	 else if (in[16:0] >= 3030 && in <= 3034) out = 2772;
	 	 	 else if (in[16:0] >= 3035 && in <= 3038) out = 2773;
	 	 	 else if (in[16:0] >= 3039 && in <= 3043) out = 2774;
	 	 	 else if (in[16:0] >= 3044 && in <= 3047) out = 2775;
	 	 	 else if (in[16:0] >= 3048 && in <= 3052) out = 2776;
	 	 	 else if (in[16:0] >= 3053 && in <= 3057) out = 2777;
	 	 	 else if (in[16:0] >= 3058 && in <= 3061) out = 2778;
	 	 	 else if (in[16:0] >= 3062 && in <= 3066) out = 2779;
	 	 	 else if (in[16:0] >= 3067 && in <= 3070) out = 2780;
	 	 	 else if (in[16:0] >= 3071 && in <= 3075) out = 2781;
	 	 	 else if (in[16:0] >= 3076 && in <= 3080) out = 2782;
	 	 	 else if (in[16:0] >= 3081 && in <= 3084) out = 2783;
	 	 	 else if (in[16:0] >= 3085 && in <= 3089) out = 2784;
	 	 	 else if (in[16:0] >= 3090 && in <= 3093) out = 2785;
	 	 	 else if (in[16:0] >= 3094 && in <= 3098) out = 2786;
	 	 	 else if (in[16:0] >= 3099 && in <= 3103) out = 2787;
	 	 	 else if (in[16:0] >= 3104 && in <= 3107) out = 2788;
	 	 	 else if (in[16:0] >= 3108 && in <= 3112) out = 2789;
	 	 	 else if (in[16:0] >= 3113 && in <= 3116) out = 2790;
	 	 	 else if (in[16:0] >= 3117 && in <= 3121) out = 2791;
	 	 	 else if (in[16:0] >= 3122 && in <= 3126) out = 2792;
	 	 	 else if (in[16:0] >= 3127 && in <= 3130) out = 2793;
	 	 	 else if (in[16:0] >= 3131 && in <= 3135) out = 2794;
	 	 	 else if (in[16:0] >= 3136 && in <= 3139) out = 2795;
	 	 	 else if (in[16:0] >= 3140 && in <= 3144) out = 2796;
	 	 	 else if (in[16:0] >= 3145 && in <= 3149) out = 2797;
	 	 	 else if (in[16:0] >= 3150 && in <= 3153) out = 2798;
	 	 	 else if (in[16:0] >= 3154 && in <= 3158) out = 2799;
	 	 	 else if (in[16:0] >= 3159 && in <= 3163) out = 2800;
	 	 	 else if (in[16:0] >= 3164 && in <= 3167) out = 2801;
	 	 	 else if (in[16:0] >= 3168 && in <= 3172) out = 2802;
	 	 	 else if (in[16:0] >= 3173 && in <= 3176) out = 2803;
	 	 	 else if (in[16:0] >= 3177 && in <= 3181) out = 2804;
	 	 	 else if (in[16:0] >= 3182 && in <= 3186) out = 2805;
	 	 	 else if (in[16:0] >= 3187 && in <= 3190) out = 2806;
	 	 	 else if (in[16:0] >= 3191 && in <= 3195) out = 2807;
	 	 	 else if (in[16:0] >= 3196 && in <= 3200) out = 2808;
	 	 	 else if (in[16:0] >= 3201 && in <= 3204) out = 2809;
	 	 	 else if (in[16:0] >= 3205 && in <= 3209) out = 2810;
	 	 	 else if (in[16:0] >= 3210 && in <= 3214) out = 2811;
	 	 	 else if (in[16:0] >= 3215 && in <= 3218) out = 2812;
	 	 	 else if (in[16:0] >= 3219 && in <= 3223) out = 2813;
	 	 	 else if (in[16:0] >= 3224 && in <= 3228) out = 2814;
	 	 	 else if (in[16:0] >= 3229 && in <= 3232) out = 2815;
	 	 	 else if (in[16:0] >= 3233 && in <= 3237) out = 2816;
	 	 	 else if (in[16:0] >= 3238 && in <= 3242) out = 2817;
	 	 	 else if (in[16:0] >= 3243 && in <= 3246) out = 2818;
	 	 	 else if (in[16:0] >= 3247 && in <= 3251) out = 2819;
	 	 	 else if (in[16:0] >= 3252 && in <= 3256) out = 2820;
	 	 	 else if (in[16:0] >= 3257 && in <= 3260) out = 2821;
	 	 	 else if (in[16:0] >= 3261 && in <= 3265) out = 2822;
	 	 	 else if (in[16:0] >= 3266 && in <= 3270) out = 2823;
	 	 	 else if (in[16:0] >= 3271 && in <= 3274) out = 2824;
	 	 	 else if (in[16:0] >= 3275 && in <= 3279) out = 2825;
	 	 	 else if (in[16:0] >= 3280 && in <= 3284) out = 2826;
	 	 	 else if (in[16:0] >= 3285 && in <= 3288) out = 2827;
	 	 	 else if (in[16:0] >= 3289 && in <= 3293) out = 2828;
	 	 	 else if (in[16:0] >= 3294 && in <= 3298) out = 2829;
	 	 	 else if (in[16:0] >= 3299 && in <= 3302) out = 2830;
	 	 	 else if (in[16:0] >= 3303 && in <= 3307) out = 2831;
	 	 	 else if (in[16:0] >= 3308 && in <= 3312) out = 2832;
	 	 	 else if (in[16:0] >= 3313 && in <= 3316) out = 2833;
	 	 	 else if (in[16:0] >= 3317 && in <= 3321) out = 2834;
	 	 	 else if (in[16:0] >= 3322 && in <= 3326) out = 2835;
	 	 	 else if (in[16:0] >= 3327 && in <= 3330) out = 2836;
	 	 	 else if (in[16:0] >= 3331 && in <= 3335) out = 2837;
	 	 	 else if (in[16:0] >= 3336 && in <= 3340) out = 2838;
	 	 	 else if (in[16:0] >= 3341 && in <= 3345) out = 2839;
	 	 	 else if (in[16:0] >= 3346 && in <= 3349) out = 2840;
	 	 	 else if (in[16:0] >= 3350 && in <= 3354) out = 2841;
	 	 	 else if (in[16:0] >= 3355 && in <= 3359) out = 2842;
	 	 	 else if (in[16:0] >= 3360 && in <= 3363) out = 2843;
	 	 	 else if (in[16:0] >= 3364 && in <= 3368) out = 2844;
	 	 	 else if (in[16:0] >= 3369 && in <= 3373) out = 2845;
	 	 	 else if (in[16:0] >= 3374 && in <= 3378) out = 2846;
	 	 	 else if (in[16:0] >= 3379 && in <= 3382) out = 2847;
	 	 	 else if (in[16:0] >= 3383 && in <= 3387) out = 2848;
	 	 	 else if (in[16:0] >= 3388 && in <= 3392) out = 2849;
	 	 	 else if (in[16:0] >= 3393 && in <= 3396) out = 2850;
	 	 	 else if (in[16:0] >= 3397 && in <= 3401) out = 2851;
	 	 	 else if (in[16:0] >= 3402 && in <= 3406) out = 2852;
	 	 	 else if (in[16:0] >= 3407 && in <= 3411) out = 2853;
	 	 	 else if (in[16:0] >= 3412 && in <= 3415) out = 2854;
	 	 	 else if (in[16:0] >= 3416 && in <= 3420) out = 2855;
	 	 	 else if (in[16:0] >= 3421 && in <= 3425) out = 2856;
	 	 	 else if (in[16:0] >= 3426 && in <= 3430) out = 2857;
	 	 	 else if (in[16:0] >= 3431 && in <= 3434) out = 2858;
	 	 	 else if (in[16:0] >= 3435 && in <= 3439) out = 2859;
	 	 	 else if (in[16:0] >= 3440 && in <= 3444) out = 2860;
	 	 	 else if (in[16:0] >= 3445 && in <= 3449) out = 2861;
	 	 	 else if (in[16:0] >= 3450 && in <= 3453) out = 2862;
	 	 	 else if (in[16:0] >= 3454 && in <= 3458) out = 2863;
	 	 	 else if (in[16:0] >= 3459 && in <= 3463) out = 2864;
	 	 	 else if (in[16:0] >= 3464 && in <= 3468) out = 2865;
	 	 	 else if (in[16:0] >= 3469 && in <= 3472) out = 2866;
	 	 	 else if (in[16:0] >= 3473 && in <= 3477) out = 2867;
	 	 	 else if (in[16:0] >= 3478 && in <= 3482) out = 2868;
	 	 	 else if (in[16:0] >= 3483 && in <= 3487) out = 2869;
	 	 	 else if (in[16:0] >= 3488 && in <= 3491) out = 2870;
	 	 	 else if (in[16:0] >= 3492 && in <= 3496) out = 2871;
	 	 	 else if (in[16:0] >= 3497 && in <= 3501) out = 2872;
	 	 	 else if (in[16:0] >= 3502 && in <= 3506) out = 2873;
	 	 	 else if (in[16:0] >= 3507 && in <= 3511) out = 2874;
	 	 	 else if (in[16:0] >= 3512 && in <= 3515) out = 2875;
	 	 	 else if (in[16:0] >= 3516 && in <= 3520) out = 2876;
	 	 	 else if (in[16:0] >= 3521 && in <= 3525) out = 2877;
	 	 	 else if (in[16:0] >= 3526 && in <= 3530) out = 2878;
	 	 	 else if (in[16:0] >= 3531 && in <= 3535) out = 2879;
	 	 	 else if (in[16:0] >= 3536 && in <= 3539) out = 2880;
	 	 	 else if (in[16:0] >= 3540 && in <= 3544) out = 2881;
	 	 	 else if (in[16:0] >= 3545 && in <= 3549) out = 2882;
	 	 	 else if (in[16:0] >= 3550 && in <= 3554) out = 2883;
	 	 	 else if (in[16:0] >= 3555 && in <= 3559) out = 2884;
	 	 	 else if (in[16:0] >= 3560 && in <= 3563) out = 2885;
	 	 	 else if (in[16:0] >= 3564 && in <= 3568) out = 2886;
	 	 	 else if (in[16:0] >= 3569 && in <= 3573) out = 2887;
	 	 	 else if (in[16:0] >= 3574 && in <= 3578) out = 2888;
	 	 	 else if (in[16:0] >= 3579 && in <= 3583) out = 2889;
	 	 	 else if (in[16:0] >= 3584 && in <= 3587) out = 2890;
	 	 	 else if (in[16:0] >= 3588 && in <= 3592) out = 2891;
	 	 	 else if (in[16:0] >= 3593 && in <= 3597) out = 2892;
	 	 	 else if (in[16:0] >= 3598 && in <= 3602) out = 2893;
	 	 	 else if (in[16:0] >= 3603 && in <= 3607) out = 2894;
	 	 	 else if (in[16:0] >= 3608 && in <= 3612) out = 2895;
	 	 	 else if (in[16:0] >= 3613 && in <= 3616) out = 2896;
	 	 	 else if (in[16:0] >= 3617 && in <= 3621) out = 2897;
	 	 	 else if (in[16:0] >= 3622 && in <= 3626) out = 2898;
	 	 	 else if (in[16:0] >= 3627 && in <= 3631) out = 2899;
	 	 	 else if (in[16:0] >= 3632 && in <= 3636) out = 2900;
	 	 	 else if (in[16:0] >= 3637 && in <= 3641) out = 2901;
	 	 	 else if (in[16:0] >= 3642 && in <= 3645) out = 2902;
	 	 	 else if (in[16:0] >= 3646 && in <= 3650) out = 2903;
	 	 	 else if (in[16:0] >= 3651 && in <= 3655) out = 2904;
	 	 	 else if (in[16:0] >= 3656 && in <= 3660) out = 2905;
	 	 	 else if (in[16:0] >= 3661 && in <= 3665) out = 2906;
	 	 	 else if (in[16:0] >= 3666 && in <= 3670) out = 2907;
	 	 	 else if (in[16:0] >= 3671 && in <= 3675) out = 2908;
	 	 	 else if (in[16:0] >= 3676 && in <= 3679) out = 2909;
	 	 	 else if (in[16:0] >= 3680 && in <= 3684) out = 2910;
	 	 	 else if (in[16:0] >= 3685 && in <= 3689) out = 2911;
	 	 	 else if (in[16:0] >= 3690 && in <= 3694) out = 2912;
	 	 	 else if (in[16:0] >= 3695 && in <= 3699) out = 2913;
	 	 	 else if (in[16:0] >= 3700 && in <= 3704) out = 2914;
	 	 	 else if (in[16:0] >= 3705 && in <= 3709) out = 2915;
	 	 	 else if (in[16:0] >= 3710 && in <= 3713) out = 2916;
	 	 	 else if (in[16:0] >= 3714 && in <= 3718) out = 2917;
	 	 	 else if (in[16:0] >= 3719 && in <= 3723) out = 2918;
	 	 	 else if (in[16:0] >= 3724 && in <= 3728) out = 2919;
	 	 	 else if (in[16:0] >= 3729 && in <= 3733) out = 2920;
	 	 	 else if (in[16:0] >= 3734 && in <= 3738) out = 2921;
	 	 	 else if (in[16:0] >= 3739 && in <= 3743) out = 2922;
	 	 	 else if (in[16:0] >= 3744 && in <= 3748) out = 2923;
	 	 	 else if (in[16:0] >= 3749 && in <= 3753) out = 2924;
	 	 	 else if (in[16:0] >= 3754 && in <= 3758) out = 2925;
	 	 	 else if (in[16:0] >= 3759 && in <= 3762) out = 2926;
	 	 	 else if (in[16:0] >= 3763 && in <= 3767) out = 2927;
	 	 	 else if (in[16:0] >= 3768 && in <= 3772) out = 2928;
	 	 	 else if (in[16:0] >= 3773 && in <= 3777) out = 2929;
	 	 	 else if (in[16:0] >= 3778 && in <= 3782) out = 2930;
	 	 	 else if (in[16:0] >= 3783 && in <= 3787) out = 2931;
	 	 	 else if (in[16:0] >= 3788 && in <= 3792) out = 2932;
	 	 	 else if (in[16:0] >= 3793 && in <= 3797) out = 2933;
	 	 	 else if (in[16:0] >= 3798 && in <= 3802) out = 2934;
	 	 	 else if (in[16:0] >= 3803 && in <= 3807) out = 2935;
	 	 	 else if (in[16:0] >= 3808 && in <= 3812) out = 2936;
	 	 	 else if (in[16:0] >= 3813 && in <= 3817) out = 2937;
	 	 	 else if (in[16:0] >= 3818 && in <= 3821) out = 2938;
	 	 	 else if (in[16:0] >= 3822 && in <= 3826) out = 2939;
	 	 	 else if (in[16:0] >= 3827 && in <= 3831) out = 2940;
	 	 	 else if (in[16:0] >= 3832 && in <= 3836) out = 2941;
	 	 	 else if (in[16:0] >= 3837 && in <= 3841) out = 2942;
	 	 	 else if (in[16:0] >= 3842 && in <= 3846) out = 2943;
	 	 	 else if (in[16:0] >= 3847 && in <= 3851) out = 2944;
	 	 	 else if (in[16:0] >= 3852 && in <= 3856) out = 2945;
	 	 	 else if (in[16:0] >= 3857 && in <= 3861) out = 2946;
	 	 	 else if (in[16:0] >= 3862 && in <= 3866) out = 2947;
	 	 	 else if (in[16:0] >= 3867 && in <= 3871) out = 2948;
	 	 	 else if (in[16:0] >= 3872 && in <= 3876) out = 2949;
	 	 	 else if (in[16:0] >= 3877 && in <= 3881) out = 2950;
	 	 	 else if (in[16:0] >= 3882 && in <= 3886) out = 2951;
	 	 	 else if (in[16:0] >= 3887 && in <= 3891) out = 2952;
	 	 	 else if (in[16:0] >= 3892 && in <= 3896) out = 2953;
	 	 	 else if (in[16:0] >= 3897 && in <= 3901) out = 2954;
	 	 	 else if (in[16:0] >= 3902 && in <= 3906) out = 2955;
	 	 	 else if (in[16:0] >= 3907 && in <= 3911) out = 2956;
	 	 	 else if (in[16:0] >= 3912 && in <= 3916) out = 2957;
	 	 	 else if (in[16:0] >= 3917 && in <= 3921) out = 2958;
	 	 	 else if (in[16:0] >= 3922 && in <= 3926) out = 2959;
	 	 	 else if (in[16:0] >= 3927 && in <= 3931) out = 2960;
	 	 	 else if (in[16:0] >= 3932 && in <= 3936) out = 2961;
	 	 	 else if (in[16:0] >= 3937 && in <= 3941) out = 2962;
	 	 	 else if (in[16:0] >= 3942 && in <= 3946) out = 2963;
	 	 	 else if (in[16:0] >= 3947 && in <= 3951) out = 2964;
	 	 	 else if (in[16:0] >= 3952 && in <= 3956) out = 2965;
	 	 	 else if (in[16:0] >= 3957 && in <= 3961) out = 2966;
	 	 	 else if (in[16:0] >= 3962 && in <= 3966) out = 2967;
	 	 	 else if (in[16:0] >= 3967 && in <= 3971) out = 2968;
	 	 	 else if (in[16:0] >= 3972 && in <= 3976) out = 2969;
	 	 	 else if (in[16:0] >= 3977 && in <= 3981) out = 2970;
	 	 	 else if (in[16:0] >= 3982 && in <= 3986) out = 2971;
	 	 	 else if (in[16:0] >= 3987 && in <= 3991) out = 2972;
	 	 	 else if (in[16:0] >= 3992 && in <= 3996) out = 2973;
	 	 	 else if (in[16:0] >= 3997 && in <= 4001) out = 2974;
	 	 	 else if (in[16:0] >= 4002 && in <= 4006) out = 2975;
	 	 	 else if (in[16:0] >= 4007 && in <= 4011) out = 2976;
	 	 	 else if (in[16:0] >= 4012 && in <= 4016) out = 2977;
	 	 	 else if (in[16:0] >= 4017 && in <= 4021) out = 2978;
	 	 	 else if (in[16:0] >= 4022 && in <= 4026) out = 2979;
	 	 	 else if (in[16:0] >= 4027 && in <= 4031) out = 2980;
	 	 	 else if (in[16:0] >= 4032 && in <= 4036) out = 2981;
	 	 	 else if (in[16:0] >= 4037 && in <= 4041) out = 2982;
	 	 	 else if (in[16:0] >= 4042 && in <= 4046) out = 2983;
	 	 	 else if (in[16:0] >= 4047 && in <= 4051) out = 2984;
	 	 	 else if (in[16:0] >= 4052 && in <= 4056) out = 2985;
	 	 	 else if (in[16:0] >= 4057 && in <= 4062) out = 2986;
	 	 	 else if (in[16:0] >= 4063 && in <= 4067) out = 2987;
	 	 	 else if (in[16:0] >= 4068 && in <= 4072) out = 2988;
	 	 	 else if (in[16:0] >= 4073 && in <= 4077) out = 2989;
	 	 	 else if (in[16:0] >= 4078 && in <= 4082) out = 2990;
	 	 	 else if (in[16:0] >= 4083 && in <= 4087) out = 2991;
	 	 	 else if (in[16:0] >= 4088 && in <= 4092) out = 2992;
	 	 	 else if (in[16:0] >= 4093 && in <= 4097) out = 2993;
	 	 	 else if (in[16:0] >= 4098 && in <= 4102) out = 2994;
	 	 	 else if (in[16:0] >= 4103 && in <= 4107) out = 2995;
	 	 	 else if (in[16:0] >= 4108 && in <= 4112) out = 2996;
	 	 	 else if (in[16:0] >= 4113 && in <= 4117) out = 2997;
	 	 	 else if (in[16:0] >= 4118 && in <= 4123) out = 2998;
	 	 	 else if (in[16:0] >= 4124 && in <= 4128) out = 2999;
	 	 	 else if (in[16:0] >= 4129 && in <= 4133) out = 3000;
	 	 	 else if (in[16:0] >= 4134 && in <= 4138) out = 3001;
	 	 	 else if (in[16:0] >= 4139 && in <= 4143) out = 3002;
	 	 	 else if (in[16:0] >= 4144 && in <= 4148) out = 3003;
	 	 	 else if (in[16:0] >= 4149 && in <= 4153) out = 3004;
	 	 	 else if (in[16:0] >= 4154 && in <= 4158) out = 3005;
	 	 	 else if (in[16:0] >= 4159 && in <= 4164) out = 3006;
	 	 	 else if (in[16:0] >= 4165 && in <= 4169) out = 3007;
	 	 	 else if (in[16:0] >= 4170 && in <= 4174) out = 3008;
	 	 	 else if (in[16:0] >= 4175 && in <= 4179) out = 3009;
	 	 	 else if (in[16:0] >= 4180 && in <= 4184) out = 3010;
	 	 	 else if (in[16:0] >= 4185 && in <= 4189) out = 3011;
	 	 	 else if (in[16:0] >= 4190 && in <= 4194) out = 3012;
	 	 	 else if (in[16:0] >= 4195 && in <= 4199) out = 3013;
	 	 	 else if (in[16:0] >= 4200 && in <= 4205) out = 3014;
	 	 	 else if (in[16:0] >= 4206 && in <= 4210) out = 3015;
	 	 	 else if (in[16:0] >= 4211 && in <= 4215) out = 3016;
	 	 	 else if (in[16:0] >= 4216 && in <= 4220) out = 3017;
	 	 	 else if (in[16:0] >= 4221 && in <= 4225) out = 3018;
	 	 	 else if (in[16:0] >= 4226 && in <= 4230) out = 3019;
	 	 	 else if (in[16:0] >= 4231 && in <= 4236) out = 3020;
	 	 	 else if (in[16:0] >= 4237 && in <= 4241) out = 3021;
	 	 	 else if (in[16:0] >= 4242 && in <= 4246) out = 3022;
	 	 	 else if (in[16:0] >= 4247 && in <= 4251) out = 3023;
	 	 	 else if (in[16:0] >= 4252 && in <= 4256) out = 3024;
	 	 	 else if (in[16:0] >= 4257 && in <= 4261) out = 3025;
	 	 	 else if (in[16:0] >= 4262 && in <= 4267) out = 3026;
	 	 	 else if (in[16:0] >= 4268 && in <= 4272) out = 3027;
	 	 	 else if (in[16:0] >= 4273 && in <= 4277) out = 3028;
	 	 	 else if (in[16:0] >= 4278 && in <= 4282) out = 3029;
	 	 	 else if (in[16:0] >= 4283 && in <= 4287) out = 3030;
	 	 	 else if (in[16:0] >= 4288 && in <= 4293) out = 3031;
	 	 	 else if (in[16:0] >= 4294 && in <= 4298) out = 3032;
	 	 	 else if (in[16:0] >= 4299 && in <= 4303) out = 3033;
	 	 	 else if (in[16:0] >= 4304 && in <= 4308) out = 3034;
	 	 	 else if (in[16:0] >= 4309 && in <= 4313) out = 3035;
	 	 	 else if (in[16:0] >= 4314 && in <= 4319) out = 3036;
	 	 	 else if (in[16:0] >= 4320 && in <= 4324) out = 3037;
	 	 	 else if (in[16:0] >= 4325 && in <= 4329) out = 3038;
	 	 	 else if (in[16:0] >= 4330 && in <= 4334) out = 3039;
	 	 	 else if (in[16:0] >= 4335 && in <= 4340) out = 3040;
	 	 	 else if (in[16:0] >= 4341 && in <= 4345) out = 3041;
	 	 	 else if (in[16:0] >= 4346 && in <= 4350) out = 3042;
	 	 	 else if (in[16:0] >= 4351 && in <= 4355) out = 3043;
	 	 	 else if (in[16:0] >= 4356 && in <= 4361) out = 3044;
	 	 	 else if (in[16:0] >= 4362 && in <= 4366) out = 3045;
	 	 	 else if (in[16:0] >= 4367 && in <= 4371) out = 3046;
	 	 	 else if (in[16:0] >= 4372 && in <= 4376) out = 3047;
	 	 	 else if (in[16:0] >= 4377 && in <= 4382) out = 3048;
	 	 	 else if (in[16:0] >= 4383 && in <= 4387) out = 3049;
	 	 	 else if (in[16:0] >= 4388 && in <= 4392) out = 3050;
	 	 	 else if (in[16:0] >= 4393 && in <= 4397) out = 3051;
	 	 	 else if (in[16:0] >= 4398 && in <= 4403) out = 3052;
	 	 	 else if (in[16:0] >= 4404 && in <= 4408) out = 3053;
	 	 	 else if (in[16:0] >= 4409 && in <= 4413) out = 3054;
	 	 	 else if (in[16:0] >= 4414 && in <= 4418) out = 3055;
	 	 	 else if (in[16:0] >= 4419 && in <= 4424) out = 3056;
	 	 	 else if (in[16:0] >= 4425 && in <= 4429) out = 3057;
	 	 	 else if (in[16:0] >= 4430 && in <= 4434) out = 3058;
	 	 	 else if (in[16:0] >= 4435 && in <= 4440) out = 3059;
	 	 	 else if (in[16:0] >= 4441 && in <= 4445) out = 3060;
	 	 	 else if (in[16:0] >= 4446 && in <= 4450) out = 3061;
	 	 	 else if (in[16:0] >= 4451 && in <= 4456) out = 3062;
	 	 	 else if (in[16:0] >= 4457 && in <= 4461) out = 3063;
	 	 	 else if (in[16:0] >= 4462 && in <= 4466) out = 3064;
	 	 	 else if (in[16:0] >= 4467 && in <= 4471) out = 3065;
	 	 	 else if (in[16:0] >= 4472 && in <= 4477) out = 3066;
	 	 	 else if (in[16:0] >= 4478 && in <= 4482) out = 3067;
	 	 	 else if (in[16:0] >= 4483 && in <= 4487) out = 3068;
	 	 	 else if (in[16:0] >= 4488 && in <= 4493) out = 3069;
	 	 	 else if (in[16:0] >= 4494 && in <= 4498) out = 3070;
	 	 	 else if (in[16:0] >= 4499 && in <= 4503) out = 3071;
	 	 	 else if (in[16:0] >= 4504 && in <= 4509) out = 3072;
	 	 	 else if (in[16:0] >= 4510 && in <= 4514) out = 3073;
	 	 	 else if (in[16:0] >= 4515 && in <= 4519) out = 3074;
	 	 	 else if (in[16:0] >= 4520 && in <= 4525) out = 3075;
	 	 	 else if (in[16:0] >= 4526 && in <= 4530) out = 3076;
	 	 	 else if (in[16:0] >= 4531 && in <= 4536) out = 3077;
	 	 	 else if (in[16:0] >= 4537 && in <= 4541) out = 3078;
	 	 	 else if (in[16:0] >= 4542 && in <= 4546) out = 3079;
	 	 	 else if (in[16:0] >= 4547 && in <= 4552) out = 3080;
	 	 	 else if (in[16:0] >= 4553 && in <= 4557) out = 3081;
	 	 	 else if (in[16:0] >= 4558 && in <= 4562) out = 3082;
	 	 	 else if (in[16:0] >= 4563 && in <= 4568) out = 3083;
	 	 	 else if (in[16:0] >= 4569 && in <= 4573) out = 3084;
	 	 	 else if (in[16:0] >= 4574 && in <= 4578) out = 3085;
	 	 	 else if (in[16:0] >= 4579 && in <= 4584) out = 3086;
	 	 	 else if (in[16:0] >= 4585 && in <= 4589) out = 3087;
	 	 	 else if (in[16:0] >= 4590 && in <= 4595) out = 3088;
	 	 	 else if (in[16:0] >= 4596 && in <= 4600) out = 3089;
	 	 	 else if (in[16:0] >= 4601 && in <= 4605) out = 3090;
	 	 	 else if (in[16:0] >= 4606 && in <= 4611) out = 3091;
	 	 	 else if (in[16:0] >= 4612 && in <= 4616) out = 3092;
	 	 	 else if (in[16:0] >= 4617 && in <= 4622) out = 3093;
	 	 	 else if (in[16:0] >= 4623 && in <= 4627) out = 3094;
	 	 	 else if (in[16:0] >= 4628 && in <= 4633) out = 3095;
	 	 	 else if (in[16:0] >= 4634 && in <= 4638) out = 3096;
	 	 	 else if (in[16:0] >= 4639 && in <= 4643) out = 3097;
	 	 	 else if (in[16:0] >= 4644 && in <= 4649) out = 3098;
	 	 	 else if (in[16:0] >= 4650 && in <= 4654) out = 3099;
	 	 	 else if (in[16:0] >= 4655 && in <= 4660) out = 3100;
	 	 	 else if (in[16:0] >= 4661 && in <= 4665) out = 3101;
	 	 	 else if (in[16:0] >= 4666 && in <= 4671) out = 3102;
	 	 	 else if (in[16:0] >= 4672 && in <= 4676) out = 3103;
	 	 	 else if (in[16:0] >= 4677 && in <= 4681) out = 3104;
	 	 	 else if (in[16:0] >= 4682 && in <= 4687) out = 3105;
	 	 	 else if (in[16:0] >= 4688 && in <= 4692) out = 3106;
	 	 	 else if (in[16:0] >= 4693 && in <= 4698) out = 3107;
	 	 	 else if (in[16:0] >= 4699 && in <= 4703) out = 3108;
	 	 	 else if (in[16:0] >= 4704 && in <= 4709) out = 3109;
	 	 	 else if (in[16:0] >= 4710 && in <= 4714) out = 3110;
	 	 	 else if (in[16:0] >= 4715 && in <= 4720) out = 3111;
	 	 	 else if (in[16:0] >= 4721 && in <= 4725) out = 3112;
	 	 	 else if (in[16:0] >= 4726 && in <= 4731) out = 3113;
	 	 	 else if (in[16:0] >= 4732 && in <= 4736) out = 3114;
	 	 	 else if (in[16:0] >= 4737 && in <= 4742) out = 3115;
	 	 	 else if (in[16:0] >= 4743 && in <= 4747) out = 3116;
	 	 	 else if (in[16:0] >= 4748 && in <= 4753) out = 3117;
	 	 	 else if (in[16:0] >= 4754 && in <= 4758) out = 3118;
	 	 	 else if (in[16:0] >= 4759 && in <= 4764) out = 3119;
	 	 	 else if (in[16:0] >= 4765 && in <= 4769) out = 3120;
	 	 	 else if (in[16:0] >= 4770 && in <= 4775) out = 3121;
	 	 	 else if (in[16:0] >= 4776 && in <= 4780) out = 3122;
	 	 	 else if (in[16:0] >= 4781 && in <= 4786) out = 3123;
	 	 	 else if (in[16:0] >= 4787 && in <= 4791) out = 3124;
	 	 	 else if (in[16:0] >= 4792 && in <= 4797) out = 3125;
	 	 	 else if (in[16:0] >= 4798 && in <= 4802) out = 3126;
	 	 	 else if (in[16:0] >= 4803 && in <= 4808) out = 3127;
	 	 	 else if (in[16:0] >= 4809 && in <= 4814) out = 3128;
	 	 	 else if (in[16:0] >= 4815 && in <= 4819) out = 3129;
	 	 	 else if (in[16:0] >= 4820 && in <= 4825) out = 3130;
	 	 	 else if (in[16:0] >= 4826 && in <= 4830) out = 3131;
	 	 	 else if (in[16:0] >= 4831 && in <= 4836) out = 3132;
	 	 	 else if (in[16:0] >= 4837 && in <= 4841) out = 3133;
	 	 	 else if (in[16:0] >= 4842 && in <= 4847) out = 3134;
	 	 	 else if (in[16:0] >= 4848 && in <= 4852) out = 3135;
	 	 	 else if (in[16:0] >= 4853 && in <= 4858) out = 3136;
	 	 	 else if (in[16:0] >= 4859 && in <= 4864) out = 3137;
	 	 	 else if (in[16:0] >= 4865 && in <= 4869) out = 3138;
	 	 	 else if (in[16:0] >= 4870 && in <= 4875) out = 3139;
	 	 	 else if (in[16:0] >= 4876 && in <= 4880) out = 3140;
	 	 	 else if (in[16:0] >= 4881 && in <= 4886) out = 3141;
	 	 	 else if (in[16:0] >= 4887 && in <= 4892) out = 3142;
	 	 	 else if (in[16:0] >= 4893 && in <= 4897) out = 3143;
	 	 	 else if (in[16:0] >= 4898 && in <= 4903) out = 3144;
	 	 	 else if (in[16:0] >= 4904 && in <= 4908) out = 3145;
	 	 	 else if (in[16:0] >= 4909 && in <= 4914) out = 3146;
	 	 	 else if (in[16:0] >= 4915 && in <= 4920) out = 3147;
	 	 	 else if (in[16:0] >= 4921 && in <= 4925) out = 3148;
	 	 	 else if (in[16:0] >= 4926 && in <= 4931) out = 3149;
	 	 	 else if (in[16:0] >= 4932 && in <= 4937) out = 3150;
	 	 	 else if (in[16:0] >= 4938 && in <= 4942) out = 3151;
	 	 	 else if (in[16:0] >= 4943 && in <= 4948) out = 3152;
	 	 	 else if (in[16:0] >= 4949 && in <= 4954) out = 3153;
	 	 	 else if (in[16:0] >= 4955 && in <= 4959) out = 3154;
	 	 	 else if (in[16:0] >= 4960 && in <= 4965) out = 3155;
	 	 	 else if (in[16:0] >= 4966 && in <= 4971) out = 3156;
	 	 	 else if (in[16:0] >= 4972 && in <= 4976) out = 3157;
	 	 	 else if (in[16:0] >= 4977 && in <= 4982) out = 3158;
	 	 	 else if (in[16:0] >= 4983 && in <= 4988) out = 3159;
	 	 	 else if (in[16:0] >= 4989 && in <= 4993) out = 3160;
	 	 	 else if (in[16:0] >= 4994 && in <= 4999) out = 3161;
	 	 	 else if (in[16:0] >= 5000 && in <= 5005) out = 3162;
	 	 	 else if (in[16:0] >= 5006 && in <= 5010) out = 3163;
	 	 	 else if (in[16:0] >= 5011 && in <= 5016) out = 3164;
	 	 	 else if (in[16:0] >= 5017 && in <= 5022) out = 3165;
	 	 	 else if (in[16:0] >= 5023 && in <= 5027) out = 3166;
	 	 	 else if (in[16:0] >= 5028 && in <= 5033) out = 3167;
	 	 	 else if (in[16:0] >= 5034 && in <= 5039) out = 3168;
	 	 	 else if (in[16:0] >= 5040 && in <= 5045) out = 3169;
	 	 	 else if (in[16:0] >= 5046 && in <= 5050) out = 3170;
	 	 	 else if (in[16:0] >= 5051 && in <= 5056) out = 3171;
	 	 	 else if (in[16:0] >= 5057 && in <= 5062) out = 3172;
	 	 	 else if (in[16:0] >= 5063 && in <= 5067) out = 3173;
	 	 	 else if (in[16:0] >= 5068 && in <= 5073) out = 3174;
	 	 	 else if (in[16:0] >= 5074 && in <= 5079) out = 3175;
	 	 	 else if (in[16:0] >= 5080 && in <= 5085) out = 3176;
	 	 	 else if (in[16:0] >= 5086 && in <= 5090) out = 3177;
	 	 	 else if (in[16:0] >= 5091 && in <= 5096) out = 3178;
	 	 	 else if (in[16:0] >= 5097 && in <= 5102) out = 3179;
	 	 	 else if (in[16:0] >= 5103 && in <= 5108) out = 3180;
	 	 	 else if (in[16:0] >= 5109 && in <= 5113) out = 3181;
	 	 	 else if (in[16:0] >= 5114 && in <= 5119) out = 3182;
	 	 	 else if (in[16:0] >= 5120 && in <= 5125) out = 3183;
	 	 	 else if (in[16:0] >= 5126 && in <= 5131) out = 3184;
	 	 	 else if (in[16:0] >= 5132 && in <= 5137) out = 3185;
	 	 	 else if (in[16:0] >= 5138 && in <= 5142) out = 3186;
	 	 	 else if (in[16:0] >= 5143 && in <= 5148) out = 3187;
	 	 	 else if (in[16:0] >= 5149 && in <= 5154) out = 3188;
	 	 	 else if (in[16:0] >= 5155 && in <= 5160) out = 3189;
	 	 	 else if (in[16:0] >= 5161 && in <= 5166) out = 3190;
	 	 	 else if (in[16:0] >= 5167 && in <= 5171) out = 3191;
	 	 	 else if (in[16:0] >= 5172 && in <= 5177) out = 3192;
	 	 	 else if (in[16:0] >= 5178 && in <= 5183) out = 3193;
	 	 	 else if (in[16:0] >= 5184 && in <= 5189) out = 3194;
	 	 	 else if (in[16:0] >= 5190 && in <= 5195) out = 3195;
	 	 	 else if (in[16:0] >= 5196 && in <= 5201) out = 3196;
	 	 	 else if (in[16:0] >= 5202 && in <= 5206) out = 3197;
	 	 	 else if (in[16:0] >= 5207 && in <= 5212) out = 3198;
	 	 	 else if (in[16:0] >= 5213 && in <= 5218) out = 3199;
	 	 	 else if (in[16:0] >= 5219 && in <= 5224) out = 3200;
	 	 	 else if (in[16:0] >= 5225 && in <= 5230) out = 3201;
	 	 	 else if (in[16:0] >= 5231 && in <= 5236) out = 3202;
	 	 	 else if (in[16:0] >= 5237 && in <= 5242) out = 3203;
	 	 	 else if (in[16:0] >= 5243 && in <= 5247) out = 3204;
	 	 	 else if (in[16:0] >= 5248 && in <= 5253) out = 3205;
	 	 	 else if (in[16:0] >= 5254 && in <= 5259) out = 3206;
	 	 	 else if (in[16:0] >= 5260 && in <= 5265) out = 3207;
	 	 	 else if (in[16:0] >= 5266 && in <= 5271) out = 3208;
	 	 	 else if (in[16:0] >= 5272 && in <= 5277) out = 3209;
	 	 	 else if (in[16:0] >= 5278 && in <= 5283) out = 3210;
	 	 	 else if (in[16:0] >= 5284 && in <= 5289) out = 3211;
	 	 	 else if (in[16:0] >= 5290 && in <= 5295) out = 3212;
	 	 	 else if (in[16:0] >= 5296 && in <= 5301) out = 3213;
	 	 	 else if (in[16:0] >= 5302 && in <= 5307) out = 3214;
	 	 	 else if (in[16:0] >= 5308 && in <= 5312) out = 3215;
	 	 	 else if (in[16:0] >= 5313 && in <= 5318) out = 3216;
	 	 	 else if (in[16:0] >= 5319 && in <= 5324) out = 3217;
	 	 	 else if (in[16:0] >= 5325 && in <= 5330) out = 3218;
	 	 	 else if (in[16:0] >= 5331 && in <= 5336) out = 3219;
	 	 	 else if (in[16:0] >= 5337 && in <= 5342) out = 3220;
	 	 	 else if (in[16:0] >= 5343 && in <= 5348) out = 3221;
	 	 	 else if (in[16:0] >= 5349 && in <= 5354) out = 3222;
	 	 	 else if (in[16:0] >= 5355 && in <= 5360) out = 3223;
	 	 	 else if (in[16:0] >= 5361 && in <= 5366) out = 3224;
	 	 	 else if (in[16:0] >= 5367 && in <= 5372) out = 3225;
	 	 	 else if (in[16:0] >= 5373 && in <= 5378) out = 3226;
	 	 	 else if (in[16:0] >= 5379 && in <= 5384) out = 3227;
	 	 	 else if (in[16:0] >= 5385 && in <= 5390) out = 3228;
	 	 	 else if (in[16:0] >= 5391 && in <= 5396) out = 3229;
	 	 	 else if (in[16:0] >= 5397 && in <= 5402) out = 3230;
	 	 	 else if (in[16:0] >= 5403 && in <= 5408) out = 3231;
	 	 	 else if (in[16:0] >= 5409 && in <= 5414) out = 3232;
	 	 	 else if (in[16:0] >= 5415 && in <= 5420) out = 3233;
	 	 	 else if (in[16:0] >= 5421 && in <= 5426) out = 3234;
	 	 	 else if (in[16:0] >= 5427 && in <= 5432) out = 3235;
	 	 	 else if (in[16:0] >= 5433 && in <= 5438) out = 3236;
	 	 	 else if (in[16:0] >= 5439 && in <= 5444) out = 3237;
	 	 	 else if (in[16:0] >= 5445 && in <= 5450) out = 3238;
	 	 	 else if (in[16:0] >= 5451 && in <= 5456) out = 3239;
	 	 	 else if (in[16:0] >= 5457 && in <= 5462) out = 3240;
	 	 	 else if (in[16:0] >= 5463 && in <= 5468) out = 3241;
	 	 	 else if (in[16:0] >= 5469 && in <= 5474) out = 3242;
	 	 	 else if (in[16:0] >= 5475 && in <= 5481) out = 3243;
	 	 	 else if (in[16:0] >= 5482 && in <= 5487) out = 3244;
	 	 	 else if (in[16:0] >= 5488 && in <= 5493) out = 3245;
	 	 	 else if (in[16:0] >= 5494 && in <= 5499) out = 3246;
	 	 	 else if (in[16:0] >= 5500 && in <= 5505) out = 3247;
	 	 	 else if (in[16:0] >= 5506 && in <= 5511) out = 3248;
	 	 	 else if (in[16:0] >= 5512 && in <= 5517) out = 3249;
	 	 	 else if (in[16:0] >= 5518 && in <= 5523) out = 3250;
	 	 	 else if (in[16:0] >= 5524 && in <= 5529) out = 3251;
	 	 	 else if (in[16:0] >= 5530 && in <= 5535) out = 3252;
	 	 	 else if (in[16:0] >= 5536 && in <= 5542) out = 3253;
	 	 	 else if (in[16:0] >= 5543 && in <= 5548) out = 3254;
	 	 	 else if (in[16:0] >= 5549 && in <= 5554) out = 3255;
	 	 	 else if (in[16:0] >= 5555 && in <= 5560) out = 3256;
	 	 	 else if (in[16:0] >= 5561 && in <= 5566) out = 3257;
	 	 	 else if (in[16:0] >= 5567 && in <= 5572) out = 3258;
	 	 	 else if (in[16:0] >= 5573 && in <= 5578) out = 3259;
	 	 	 else if (in[16:0] >= 5579 && in <= 5585) out = 3260;
	 	 	 else if (in[16:0] >= 5586 && in <= 5591) out = 3261;
	 	 	 else if (in[16:0] >= 5592 && in <= 5597) out = 3262;
	 	 	 else if (in[16:0] >= 5598 && in <= 5603) out = 3263;
	 	 	 else if (in[16:0] >= 5604 && in <= 5609) out = 3264;
	 	 	 else if (in[16:0] >= 5610 && in <= 5616) out = 3265;
	 	 	 else if (in[16:0] >= 5617 && in <= 5622) out = 3266;
	 	 	 else if (in[16:0] >= 5623 && in <= 5628) out = 3267;
	 	 	 else if (in[16:0] >= 5629 && in <= 5634) out = 3268;
	 	 	 else if (in[16:0] >= 5635 && in <= 5640) out = 3269;
	 	 	 else if (in[16:0] >= 5641 && in <= 5647) out = 3270;
	 	 	 else if (in[16:0] >= 5648 && in <= 5653) out = 3271;
	 	 	 else if (in[16:0] >= 5654 && in <= 5659) out = 3272;
	 	 	 else if (in[16:0] >= 5660 && in <= 5665) out = 3273;
	 	 	 else if (in[16:0] >= 5666 && in <= 5672) out = 3274;
	 	 	 else if (in[16:0] >= 5673 && in <= 5678) out = 3275;
	 	 	 else if (in[16:0] >= 5679 && in <= 5684) out = 3276;
	 	 	 else if (in[16:0] >= 5685 && in <= 5690) out = 3277;
	 	 	 else if (in[16:0] >= 5691 && in <= 5697) out = 3278;
	 	 	 else if (in[16:0] >= 5698 && in <= 5703) out = 3279;
	 	 	 else if (in[16:0] >= 5704 && in <= 5709) out = 3280;
	 	 	 else if (in[16:0] >= 5710 && in <= 5715) out = 3281;
	 	 	 else if (in[16:0] >= 5716 && in <= 5722) out = 3282;
	 	 	 else if (in[16:0] >= 5723 && in <= 5728) out = 3283;
	 	 	 else if (in[16:0] >= 5729 && in <= 5734) out = 3284;
	 	 	 else if (in[16:0] >= 5735 && in <= 5741) out = 3285;
	 	 	 else if (in[16:0] >= 5742 && in <= 5747) out = 3286;
	 	 	 else if (in[16:0] >= 5748 && in <= 5753) out = 3287;
	 	 	 else if (in[16:0] >= 5754 && in <= 5760) out = 3288;
	 	 	 else if (in[16:0] >= 5761 && in <= 5766) out = 3289;
	 	 	 else if (in[16:0] >= 5767 && in <= 5772) out = 3290;
	 	 	 else if (in[16:0] >= 5773 && in <= 5779) out = 3291;
	 	 	 else if (in[16:0] >= 5780 && in <= 5785) out = 3292;
	 	 	 else if (in[16:0] >= 5786 && in <= 5791) out = 3293;
	 	 	 else if (in[16:0] >= 5792 && in <= 5798) out = 3294;
	 	 	 else if (in[16:0] >= 5799 && in <= 5804) out = 3295;
	 	 	 else if (in[16:0] >= 5805 && in <= 5810) out = 3296;
	 	 	 else if (in[16:0] >= 5811 && in <= 5817) out = 3297;
	 	 	 else if (in[16:0] >= 5818 && in <= 5823) out = 3298;
	 	 	 else if (in[16:0] >= 5824 && in <= 5829) out = 3299;
	 	 	 else if (in[16:0] >= 5830 && in <= 5836) out = 3300;
	 	 	 else if (in[16:0] >= 5837 && in <= 5842) out = 3301;
	 	 	 else if (in[16:0] >= 5843 && in <= 5849) out = 3302;
	 	 	 else if (in[16:0] >= 5850 && in <= 5855) out = 3303;
	 	 	 else if (in[16:0] >= 5856 && in <= 5862) out = 3304;
	 	 	 else if (in[16:0] >= 5863 && in <= 5868) out = 3305;
	 	 	 else if (in[16:0] >= 5869 && in <= 5874) out = 3306;
	 	 	 else if (in[16:0] >= 5875 && in <= 5881) out = 3307;
	 	 	 else if (in[16:0] >= 5882 && in <= 5887) out = 3308;
	 	 	 else if (in[16:0] >= 5888 && in <= 5894) out = 3309;
	 	 	 else if (in[16:0] >= 5895 && in <= 5900) out = 3310;
	 	 	 else if (in[16:0] >= 5901 && in <= 5907) out = 3311;
	 	 	 else if (in[16:0] >= 5908 && in <= 5913) out = 3312;
	 	 	 else if (in[16:0] >= 5914 && in <= 5920) out = 3313;
	 	 	 else if (in[16:0] >= 5921 && in <= 5926) out = 3314;
	 	 	 else if (in[16:0] >= 5927 && in <= 5933) out = 3315;
	 	 	 else if (in[16:0] >= 5934 && in <= 5939) out = 3316;
	 	 	 else if (in[16:0] >= 5940 && in <= 5946) out = 3317;
	 	 	 else if (in[16:0] >= 5947 && in <= 5952) out = 3318;
	 	 	 else if (in[16:0] >= 5953 && in <= 5959) out = 3319;
	 	 	 else if (in[16:0] >= 5960 && in <= 5965) out = 3320;
	 	 	 else if (in[16:0] >= 5966 && in <= 5972) out = 3321;
	 	 	 else if (in[16:0] >= 5973 && in <= 5978) out = 3322;
	 	 	 else if (in[16:0] >= 5979 && in <= 5985) out = 3323;
	 	 	 else if (in[16:0] >= 5986 && in <= 5991) out = 3324;
	 	 	 else if (in[16:0] >= 5992 && in <= 5998) out = 3325;
	 	 	 else if (in[16:0] >= 5999 && in <= 6004) out = 3326;
	 	 	 else if (in[16:0] >= 6005 && in <= 6011) out = 3327;
	 	 	 else if (in[16:0] >= 6012 && in <= 6018) out = 3328;
	 	 	 else if (in[16:0] >= 6019 && in <= 6024) out = 3329;
	 	 	 else if (in[16:0] >= 6025 && in <= 6031) out = 3330;
	 	 	 else if (in[16:0] >= 6032 && in <= 6037) out = 3331;
	 	 	 else if (in[16:0] >= 6038 && in <= 6044) out = 3332;
	 	 	 else if (in[16:0] >= 6045 && in <= 6050) out = 3333;
	 	 	 else if (in[16:0] >= 6051 && in <= 6057) out = 3334;
	 	 	 else if (in[16:0] >= 6058 && in <= 6064) out = 3335;
	 	 	 else if (in[16:0] >= 6065 && in <= 6070) out = 3336;
	 	 	 else if (in[16:0] >= 6071 && in <= 6077) out = 3337;
	 	 	 else if (in[16:0] >= 6078 && in <= 6084) out = 3338;
	 	 	 else if (in[16:0] >= 6085 && in <= 6090) out = 3339;
	 	 	 else if (in[16:0] >= 6091 && in <= 6097) out = 3340;
	 	 	 else if (in[16:0] >= 6098 && in <= 6104) out = 3341;
	 	 	 else if (in[16:0] >= 6105 && in <= 6110) out = 3342;
	 	 	 else if (in[16:0] >= 6111 && in <= 6117) out = 3343;
	 	 	 else if (in[16:0] >= 6118 && in <= 6124) out = 3344;
	 	 	 else if (in[16:0] >= 6125 && in <= 6130) out = 3345;
	 	 	 else if (in[16:0] >= 6131 && in <= 6137) out = 3346;
	 	 	 else if (in[16:0] >= 6138 && in <= 6144) out = 3347;
	 	 	 else if (in[16:0] >= 6145 && in <= 6150) out = 3348;
	 	 	 else if (in[16:0] >= 6151 && in <= 6157) out = 3349;
	 	 	 else if (in[16:0] >= 6158 && in <= 6164) out = 3350;
	 	 	 else if (in[16:0] >= 6165 && in <= 6171) out = 3351;
	 	 	 else if (in[16:0] >= 6172 && in <= 6177) out = 3352;
	 	 	 else if (in[16:0] >= 6178 && in <= 6184) out = 3353;
	 	 	 else if (in[16:0] >= 6185 && in <= 6191) out = 3354;
	 	 	 else if (in[16:0] >= 6192 && in <= 6198) out = 3355;
	 	 	 else if (in[16:0] >= 6199 && in <= 6204) out = 3356;
	 	 	 else if (in[16:0] >= 6205 && in <= 6211) out = 3357;
	 	 	 else if (in[16:0] >= 6212 && in <= 6218) out = 3358;
	 	 	 else if (in[16:0] >= 6219 && in <= 6225) out = 3359;
	 	 	 else if (in[16:0] >= 6226 && in <= 6232) out = 3360;
	 	 	 else if (in[16:0] >= 6233 && in <= 6238) out = 3361;
	 	 	 else if (in[16:0] >= 6239 && in <= 6245) out = 3362;
	 	 	 else if (in[16:0] >= 6246 && in <= 6252) out = 3363;
	 	 	 else if (in[16:0] >= 6253 && in <= 6259) out = 3364;
	 	 	 else if (in[16:0] >= 6260 && in <= 6266) out = 3365;
	 	 	 else if (in[16:0] >= 6267 && in <= 6272) out = 3366;
	 	 	 else if (in[16:0] >= 6273 && in <= 6279) out = 3367;
	 	 	 else if (in[16:0] >= 6280 && in <= 6286) out = 3368;
	 	 	 else if (in[16:0] >= 6287 && in <= 6293) out = 3369;
	 	 	 else if (in[16:0] >= 6294 && in <= 6300) out = 3370;
	 	 	 else if (in[16:0] >= 6301 && in <= 6307) out = 3371;
	 	 	 else if (in[16:0] >= 6308 && in <= 6314) out = 3372;
	 	 	 else if (in[16:0] >= 6315 && in <= 6321) out = 3373;
	 	 	 else if (in[16:0] >= 6322 && in <= 6327) out = 3374;
	 	 	 else if (in[16:0] >= 6328 && in <= 6334) out = 3375;
	 	 	 else if (in[16:0] >= 6335 && in <= 6341) out = 3376;
	 	 	 else if (in[16:0] >= 6342 && in <= 6348) out = 3377;
	 	 	 else if (in[16:0] >= 6349 && in <= 6355) out = 3378;
	 	 	 else if (in[16:0] >= 6356 && in <= 6362) out = 3379;
	 	 	 else if (in[16:0] >= 6363 && in <= 6369) out = 3380;
	 	 	 else if (in[16:0] >= 6370 && in <= 6376) out = 3381;
	 	 	 else if (in[16:0] >= 6377 && in <= 6383) out = 3382;
	 	 	 else if (in[16:0] >= 6384 && in <= 6390) out = 3383;
	 	 	 else if (in[16:0] >= 6391 && in <= 6397) out = 3384;
	 	 	 else if (in[16:0] >= 6398 && in <= 6404) out = 3385;
	 	 	 else if (in[16:0] >= 6405 && in <= 6411) out = 3386;
	 	 	 else if (in[16:0] >= 6412 && in <= 6418) out = 3387;
	 	 	 else if (in[16:0] >= 6419 && in <= 6425) out = 3388;
	 	 	 else if (in[16:0] >= 6426 && in <= 6432) out = 3389;
	 	 	 else if (in[16:0] >= 6433 && in <= 6439) out = 3390;
	 	 	 else if (in[16:0] >= 6440 && in <= 6446) out = 3391;
	 	 	 else if (in[16:0] >= 6447 && in <= 6453) out = 3392;
	 	 	 else if (in[16:0] >= 6454 && in <= 6460) out = 3393;
	 	 	 else if (in[16:0] >= 6461 && in <= 6467) out = 3394;
	 	 	 else if (in[16:0] >= 6468 && in <= 6474) out = 3395;
	 	 	 else if (in[16:0] >= 6475 && in <= 6481) out = 3396;
	 	 	 else if (in[16:0] >= 6482 && in <= 6488) out = 3397;
	 	 	 else if (in[16:0] >= 6489 && in <= 6495) out = 3398;
	 	 	 else if (in[16:0] >= 6496 && in <= 6502) out = 3399;
	 	 	 else if (in[16:0] >= 6503 && in <= 6509) out = 3400;
	 	 	 else if (in[16:0] >= 6510 && in <= 6517) out = 3401;
	 	 	 else if (in[16:0] >= 6518 && in <= 6524) out = 3402;
	 	 	 else if (in[16:0] >= 6525 && in <= 6531) out = 3403;
	 	 	 else if (in[16:0] >= 6532 && in <= 6538) out = 3404;
	 	 	 else if (in[16:0] >= 6539 && in <= 6545) out = 3405;
	 	 	 else if (in[16:0] >= 6546 && in <= 6552) out = 3406;
	 	 	 else if (in[16:0] >= 6553 && in <= 6559) out = 3407;
	 	 	 else if (in[16:0] >= 6560 && in <= 6567) out = 3408;
	 	 	 else if (in[16:0] >= 6568 && in <= 6574) out = 3409;
	 	 	 else if (in[16:0] >= 6575 && in <= 6581) out = 3410;
	 	 	 else if (in[16:0] >= 6582 && in <= 6588) out = 3411;
	 	 	 else if (in[16:0] >= 6589 && in <= 6595) out = 3412;
	 	 	 else if (in[16:0] >= 6596 && in <= 6603) out = 3413;
	 	 	 else if (in[16:0] >= 6604 && in <= 6610) out = 3414;
	 	 	 else if (in[16:0] >= 6611 && in <= 6617) out = 3415;
	 	 	 else if (in[16:0] >= 6618 && in <= 6624) out = 3416;
	 	 	 else if (in[16:0] >= 6625 && in <= 6631) out = 3417;
	 	 	 else if (in[16:0] >= 6632 && in <= 6639) out = 3418;
	 	 	 else if (in[16:0] >= 6640 && in <= 6646) out = 3419;
	 	 	 else if (in[16:0] >= 6647 && in <= 6653) out = 3420;
	 	 	 else if (in[16:0] >= 6654 && in <= 6661) out = 3421;
	 	 	 else if (in[16:0] >= 6662 && in <= 6668) out = 3422;
	 	 	 else if (in[16:0] >= 6669 && in <= 6675) out = 3423;
	 	 	 else if (in[16:0] >= 6676 && in <= 6682) out = 3424;
	 	 	 else if (in[16:0] >= 6683 && in <= 6690) out = 3425;
	 	 	 else if (in[16:0] >= 6691 && in <= 6697) out = 3426;
	 	 	 else if (in[16:0] >= 6698 && in <= 6704) out = 3427;
	 	 	 else if (in[16:0] >= 6705 && in <= 6712) out = 3428;
	 	 	 else if (in[16:0] >= 6713 && in <= 6719) out = 3429;
	 	 	 else if (in[16:0] >= 6720 && in <= 6726) out = 3430;
	 	 	 else if (in[16:0] >= 6727 && in <= 6734) out = 3431;
	 	 	 else if (in[16:0] >= 6735 && in <= 6741) out = 3432;
	 	 	 else if (in[16:0] >= 6742 && in <= 6749) out = 3433;
	 	 	 else if (in[16:0] >= 6750 && in <= 6756) out = 3434;
	 	 	 else if (in[16:0] >= 6757 && in <= 6763) out = 3435;
	 	 	 else if (in[16:0] >= 6764 && in <= 6771) out = 3436;
	 	 	 else if (in[16:0] >= 6772 && in <= 6778) out = 3437;
	 	 	 else if (in[16:0] >= 6779 && in <= 6786) out = 3438;
	 	 	 else if (in[16:0] >= 6787 && in <= 6793) out = 3439;
	 	 	 else if (in[16:0] >= 6794 && in <= 6801) out = 3440;
	 	 	 else if (in[16:0] >= 6802 && in <= 6808) out = 3441;
	 	 	 else if (in[16:0] >= 6809 && in <= 6815) out = 3442;
	 	 	 else if (in[16:0] >= 6816 && in <= 6823) out = 3443;
	 	 	 else if (in[16:0] >= 6824 && in <= 6830) out = 3444;
	 	 	 else if (in[16:0] >= 6831 && in <= 6838) out = 3445;
	 	 	 else if (in[16:0] >= 6839 && in <= 6845) out = 3446;
	 	 	 else if (in[16:0] >= 6846 && in <= 6853) out = 3447;
	 	 	 else if (in[16:0] >= 6854 && in <= 6860) out = 3448;
	 	 	 else if (in[16:0] >= 6861 && in <= 6868) out = 3449;
	 	 	 else if (in[16:0] >= 6869 && in <= 6876) out = 3450;
	 	 	 else if (in[16:0] >= 6877 && in <= 6883) out = 3451;
	 	 	 else if (in[16:0] >= 6884 && in <= 6891) out = 3452;
	 	 	 else if (in[16:0] >= 6892 && in <= 6898) out = 3453;
	 	 	 else if (in[16:0] >= 6899 && in <= 6906) out = 3454;
	 	 	 else if (in[16:0] >= 6907 && in <= 6913) out = 3455;
	 	 	 else if (in[16:0] >= 6914 && in <= 6921) out = 3456;
	 	 	 else if (in[16:0] >= 6922 && in <= 6929) out = 3457;
	 	 	 else if (in[16:0] >= 6930 && in <= 6936) out = 3458;
	 	 	 else if (in[16:0] >= 6937 && in <= 6944) out = 3459;
	 	 	 else if (in[16:0] >= 6945 && in <= 6951) out = 3460;
	 	 	 else if (in[16:0] >= 6952 && in <= 6959) out = 3461;
	 	 	 else if (in[16:0] >= 6960 && in <= 6967) out = 3462;
	 	 	 else if (in[16:0] >= 6968 && in <= 6974) out = 3463;
	 	 	 else if (in[16:0] >= 6975 && in <= 6982) out = 3464;
	 	 	 else if (in[16:0] >= 6983 && in <= 6990) out = 3465;
	 	 	 else if (in[16:0] >= 6991 && in <= 6998) out = 3466;
	 	 	 else if (in[16:0] >= 6999 && in <= 7005) out = 3467;
	 	 	 else if (in[16:0] >= 7006 && in <= 7013) out = 3468;
	 	 	 else if (in[16:0] >= 7014 && in <= 7021) out = 3469;
	 	 	 else if (in[16:0] >= 7022 && in <= 7028) out = 3470;
	 	 	 else if (in[16:0] >= 7029 && in <= 7036) out = 3471;
	 	 	 else if (in[16:0] >= 7037 && in <= 7044) out = 3472;
	 	 	 else if (in[16:0] >= 7045 && in <= 7052) out = 3473;
	 	 	 else if (in[16:0] >= 7053 && in <= 7059) out = 3474;
	 	 	 else if (in[16:0] >= 7060 && in <= 7067) out = 3475;
	 	 	 else if (in[16:0] >= 7068 && in <= 7075) out = 3476;
	 	 	 else if (in[16:0] >= 7076 && in <= 7083) out = 3477;
	 	 	 else if (in[16:0] >= 7084 && in <= 7091) out = 3478;
	 	 	 else if (in[16:0] >= 7092 && in <= 7099) out = 3479;
	 	 	 else if (in[16:0] >= 7100 && in <= 7106) out = 3480;
	 	 	 else if (in[16:0] >= 7107 && in <= 7114) out = 3481;
	 	 	 else if (in[16:0] >= 7115 && in <= 7122) out = 3482;
	 	 	 else if (in[16:0] >= 7123 && in <= 7130) out = 3483;
	 	 	 else if (in[16:0] >= 7131 && in <= 7138) out = 3484;
	 	 	 else if (in[16:0] >= 7139 && in <= 7146) out = 3485;
	 	 	 else if (in[16:0] >= 7147 && in <= 7154) out = 3486;
	 	 	 else if (in[16:0] >= 7155 && in <= 7162) out = 3487;
	 	 	 else if (in[16:0] >= 7163 && in <= 7170) out = 3488;
	 	 	 else if (in[16:0] >= 7171 && in <= 7177) out = 3489;
	 	 	 else if (in[16:0] >= 7178 && in <= 7185) out = 3490;
	 	 	 else if (in[16:0] >= 7186 && in <= 7193) out = 3491;
	 	 	 else if (in[16:0] >= 7194 && in <= 7201) out = 3492;
	 	 	 else if (in[16:0] >= 7202 && in <= 7209) out = 3493;
	 	 	 else if (in[16:0] >= 7210 && in <= 7217) out = 3494;
	 	 	 else if (in[16:0] >= 7218 && in <= 7225) out = 3495;
	 	 	 else if (in[16:0] >= 7226 && in <= 7233) out = 3496;
	 	 	 else if (in[16:0] >= 7234 && in <= 7241) out = 3497;
	 	 	 else if (in[16:0] >= 7242 && in <= 7249) out = 3498;
	 	 	 else if (in[16:0] >= 7250 && in <= 7257) out = 3499;
	 	 	 else if (in[16:0] >= 7258 && in <= 7265) out = 3500;
	 	 	 else if (in[16:0] >= 7266 && in <= 7274) out = 3501;
	 	 	 else if (in[16:0] >= 7275 && in <= 7282) out = 3502;
	 	 	 else if (in[16:0] >= 7283 && in <= 7290) out = 3503;
	 	 	 else if (in[16:0] >= 7291 && in <= 7298) out = 3504;
	 	 	 else if (in[16:0] >= 7299 && in <= 7306) out = 3505;
	 	 	 else if (in[16:0] >= 7307 && in <= 7314) out = 3506;
	 	 	 else if (in[16:0] >= 7315 && in <= 7322) out = 3507;
	 	 	 else if (in[16:0] >= 7323 && in <= 7330) out = 3508;
	 	 	 else if (in[16:0] >= 7331 && in <= 7339) out = 3509;
	 	 	 else if (in[16:0] >= 7340 && in <= 7347) out = 3510;
	 	 	 else if (in[16:0] >= 7348 && in <= 7355) out = 3511;
	 	 	 else if (in[16:0] >= 7356 && in <= 7363) out = 3512;
	 	 	 else if (in[16:0] >= 7364 && in <= 7371) out = 3513;
	 	 	 else if (in[16:0] >= 7372 && in <= 7380) out = 3514;
	 	 	 else if (in[16:0] >= 7381 && in <= 7388) out = 3515;
	 	 	 else if (in[16:0] >= 7389 && in <= 7396) out = 3516;
	 	 	 else if (in[16:0] >= 7397 && in <= 7404) out = 3517;
	 	 	 else if (in[16:0] >= 7405 && in <= 7413) out = 3518;
	 	 	 else if (in[16:0] >= 7414 && in <= 7421) out = 3519;
	 	 	 else if (in[16:0] >= 7422 && in <= 7429) out = 3520;
	 	 	 else if (in[16:0] >= 7430 && in <= 7437) out = 3521;
	 	 	 else if (in[16:0] >= 7438 && in <= 7446) out = 3522;
	 	 	 else if (in[16:0] >= 7447 && in <= 7454) out = 3523;
	 	 	 else if (in[16:0] >= 7455 && in <= 7462) out = 3524;
	 	 	 else if (in[16:0] >= 7463 && in <= 7471) out = 3525;
	 	 	 else if (in[16:0] >= 7472 && in <= 7479) out = 3526;
	 	 	 else if (in[16:0] >= 7480 && in <= 7488) out = 3527;
	 	 	 else if (in[16:0] >= 7489 && in <= 7496) out = 3528;
	 	 	 else if (in[16:0] >= 7497 && in <= 7504) out = 3529;
	 	 	 else if (in[16:0] >= 7505 && in <= 7513) out = 3530;
	 	 	 else if (in[16:0] >= 7514 && in <= 7521) out = 3531;
	 	 	 else if (in[16:0] >= 7522 && in <= 7530) out = 3532;
	 	 	 else if (in[16:0] >= 7531 && in <= 7538) out = 3533;
	 	 	 else if (in[16:0] >= 7539 && in <= 7547) out = 3534;
	 	 	 else if (in[16:0] >= 7548 && in <= 7555) out = 3535;
	 	 	 else if (in[16:0] >= 7556 && in <= 7563) out = 3536;
	 	 	 else if (in[16:0] >= 7564 && in <= 7572) out = 3537;
	 	 	 else if (in[16:0] >= 7573 && in <= 7581) out = 3538;
	 	 	 else if (in[16:0] >= 7582 && in <= 7589) out = 3539;
	 	 	 else if (in[16:0] >= 7590 && in <= 7598) out = 3540;
	 	 	 else if (in[16:0] >= 7599 && in <= 7606) out = 3541;
	 	 	 else if (in[16:0] >= 7607 && in <= 7615) out = 3542;
	 	 	 else if (in[16:0] >= 7616 && in <= 7623) out = 3543;
	 	 	 else if (in[16:0] >= 7624 && in <= 7632) out = 3544;
	 	 	 else if (in[16:0] >= 7633 && in <= 7640) out = 3545;
	 	 	 else if (in[16:0] >= 7641 && in <= 7649) out = 3546;
	 	 	 else if (in[16:0] >= 7650 && in <= 7658) out = 3547;
	 	 	 else if (in[16:0] >= 7659 && in <= 7666) out = 3548;
	 	 	 else if (in[16:0] >= 7667 && in <= 7675) out = 3549;
	 	 	 else if (in[16:0] >= 7676 && in <= 7684) out = 3550;
	 	 	 else if (in[16:0] >= 7685 && in <= 7692) out = 3551;
	 	 	 else if (in[16:0] >= 7693 && in <= 7701) out = 3552;
	 	 	 else if (in[16:0] >= 7702 && in <= 7710) out = 3553;
	 	 	 else if (in[16:0] >= 7711 && in <= 7719) out = 3554;
	 	 	 else if (in[16:0] >= 7720 && in <= 7727) out = 3555;
	 	 	 else if (in[16:0] >= 7728 && in <= 7736) out = 3556;
	 	 	 else if (in[16:0] >= 7737 && in <= 7745) out = 3557;
	 	 	 else if (in[16:0] >= 7746 && in <= 7754) out = 3558;
	 	 	 else if (in[16:0] >= 7755 && in <= 7762) out = 3559;
	 	 	 else if (in[16:0] >= 7763 && in <= 7771) out = 3560;
	 	 	 else if (in[16:0] >= 7772 && in <= 7780) out = 3561;
	 	 	 else if (in[16:0] >= 7781 && in <= 7789) out = 3562;
	 	 	 else if (in[16:0] >= 7790 && in <= 7798) out = 3563;
	 	 	 else if (in[16:0] >= 7799 && in <= 7807) out = 3564;
	 	 	 else if (in[16:0] >= 7808 && in <= 7816) out = 3565;
	 	 	 else if (in[16:0] >= 7817 && in <= 7824) out = 3566;
	 	 	 else if (in[16:0] >= 7825 && in <= 7833) out = 3567;
	 	 	 else if (in[16:0] >= 7834 && in <= 7842) out = 3568;
	 	 	 else if (in[16:0] >= 7843 && in <= 7851) out = 3569;
	 	 	 else if (in[16:0] >= 7852 && in <= 7860) out = 3570;
	 	 	 else if (in[16:0] >= 7861 && in <= 7869) out = 3571;
	 	 	 else if (in[16:0] >= 7870 && in <= 7878) out = 3572;
	 	 	 else if (in[16:0] >= 7879 && in <= 7887) out = 3573;
	 	 	 else if (in[16:0] >= 7888 && in <= 7896) out = 3574;
	 	 	 else if (in[16:0] >= 7897 && in <= 7905) out = 3575;
	 	 	 else if (in[16:0] >= 7906 && in <= 7914) out = 3576;
	 	 	 else if (in[16:0] >= 7915 && in <= 7923) out = 3577;
	 	 	 else if (in[16:0] >= 7924 && in <= 7932) out = 3578;
	 	 	 else if (in[16:0] >= 7933 && in <= 7941) out = 3579;
	 	 	 else if (in[16:0] >= 7942 && in <= 7951) out = 3580;
	 	 	 else if (in[16:0] >= 7952 && in <= 7960) out = 3581;
	 	 	 else if (in[16:0] >= 7961 && in <= 7969) out = 3582;
	 	 	 else if (in[16:0] >= 7970 && in <= 7978) out = 3583;
	 	 	 else if (in[16:0] >= 7979 && in <= 7987) out = 3584;
	 	 	 else if (in[16:0] >= 7988 && in <= 7996) out = 3585;
	 	 	 else if (in[16:0] >= 7997 && in <= 8006) out = 3586;
	 	 	 else if (in[16:0] >= 8007 && in <= 8015) out = 3587;
	 	 	 else if (in[16:0] >= 8016 && in <= 8024) out = 3588;
	 	 	 else if (in[16:0] >= 8025 && in <= 8033) out = 3589;
	 	 	 else if (in[16:0] >= 8034 && in <= 8042) out = 3590;
	 	 	 else if (in[16:0] >= 8043 && in <= 8052) out = 3591;
	 	 	 else if (in[16:0] >= 8053 && in <= 8061) out = 3592;
	 	 	 else if (in[16:0] >= 8062 && in <= 8070) out = 3593;
	 	 	 else if (in[16:0] >= 8071 && in <= 8080) out = 3594;
	 	 	 else if (in[16:0] >= 8081 && in <= 8089) out = 3595;
	 	 	 else if (in[16:0] >= 8090 && in <= 8098) out = 3596;
	 	 	 else if (in[16:0] >= 8099 && in <= 8108) out = 3597;
	 	 	 else if (in[16:0] >= 8109 && in <= 8117) out = 3598;
	 	 	 else if (in[16:0] >= 8118 && in <= 8127) out = 3599;
	 	 	 else if (in[16:0] >= 8128 && in <= 8136) out = 3600;
	 	 	 else if (in[16:0] >= 8137 && in <= 8145) out = 3601;
	 	 	 else if (in[16:0] >= 8146 && in <= 8155) out = 3602;
	 	 	 else if (in[16:0] >= 8156 && in <= 8164) out = 3603;
	 	 	 else if (in[16:0] >= 8165 && in <= 8174) out = 3604;
	 	 	 else if (in[16:0] >= 8175 && in <= 8183) out = 3605;
	 	 	 else if (in[16:0] >= 8184 && in <= 8193) out = 3606;
	 	 	 else if (in[16:0] >= 8194 && in <= 8202) out = 3607;
	 	 	 else if (in[16:0] >= 8203 && in <= 8212) out = 3608;
	 	 	 else if (in[16:0] >= 8213 && in <= 8221) out = 3609;
	 	 	 else if (in[16:0] >= 8222 && in <= 8231) out = 3610;
	 	 	 else if (in[16:0] >= 8232 && in <= 8241) out = 3611;
	 	 	 else if (in[16:0] >= 8242 && in <= 8250) out = 3612;
	 	 	 else if (in[16:0] >= 8251 && in <= 8260) out = 3613;
	 	 	 else if (in[16:0] >= 8261 && in <= 8270) out = 3614;
	 	 	 else if (in[16:0] >= 8271 && in <= 8279) out = 3615;
	 	 	 else if (in[16:0] >= 8280 && in <= 8289) out = 3616;
	 	 	 else if (in[16:0] >= 8290 && in <= 8299) out = 3617;
	 	 	 else if (in[16:0] >= 8300 && in <= 8308) out = 3618;
	 	 	 else if (in[16:0] >= 8309 && in <= 8318) out = 3619;
	 	 	 else if (in[16:0] >= 8319 && in <= 8328) out = 3620;
	 	 	 else if (in[16:0] >= 8329 && in <= 8338) out = 3621;
	 	 	 else if (in[16:0] >= 8339 && in <= 8347) out = 3622;
	 	 	 else if (in[16:0] >= 8348 && in <= 8357) out = 3623;
	 	 	 else if (in[16:0] >= 8358 && in <= 8367) out = 3624;
	 	 	 else if (in[16:0] >= 8368 && in <= 8377) out = 3625;
	 	 	 else if (in[16:0] >= 8378 && in <= 8387) out = 3626;
	 	 	 else if (in[16:0] >= 8388 && in <= 8397) out = 3627;
	 	 	 else if (in[16:0] >= 8398 && in <= 8407) out = 3628;
	 	 	 else if (in[16:0] >= 8408 && in <= 8417) out = 3629;
	 	 	 else if (in[16:0] >= 8418 && in <= 8427) out = 3630;
	 	 	 else if (in[16:0] >= 8428 && in <= 8436) out = 3631;
	 	 	 else if (in[16:0] >= 8437 && in <= 8446) out = 3632;
	 	 	 else if (in[16:0] >= 8447 && in <= 8456) out = 3633;
	 	 	 else if (in[16:0] >= 8457 && in <= 8466) out = 3634;
	 	 	 else if (in[16:0] >= 8467 && in <= 8477) out = 3635;
	 	 	 else if (in[16:0] >= 8478 && in <= 8487) out = 3636;
	 	 	 else if (in[16:0] >= 8488 && in <= 8497) out = 3637;
	 	 	 else if (in[16:0] >= 8498 && in <= 8507) out = 3638;
	 	 	 else if (in[16:0] >= 8508 && in <= 8517) out = 3639;
	 	 	 else if (in[16:0] >= 8518 && in <= 8527) out = 3640;
	 	 	 else if (in[16:0] >= 8528 && in <= 8537) out = 3641;
	 	 	 else if (in[16:0] >= 8538 && in <= 8547) out = 3642;
	 	 	 else if (in[16:0] >= 8548 && in <= 8558) out = 3643;
	 	 	 else if (in[16:0] >= 8559 && in <= 8568) out = 3644;
	 	 	 else if (in[16:0] >= 8569 && in <= 8578) out = 3645;
	 	 	 else if (in[16:0] >= 8579 && in <= 8588) out = 3646;
	 	 	 else if (in[16:0] >= 8589 && in <= 8599) out = 3647;
	 	 	 else if (in[16:0] >= 8600 && in <= 8609) out = 3648;
	 	 	 else if (in[16:0] >= 8610 && in <= 8619) out = 3649;
	 	 	 else if (in[16:0] >= 8620 && in <= 8629) out = 3650;
	 	 	 else if (in[16:0] >= 8630 && in <= 8640) out = 3651;
	 	 	 else if (in[16:0] >= 8641 && in <= 8650) out = 3652;
	 	 	 else if (in[16:0] >= 8651 && in <= 8661) out = 3653;
	 	 	 else if (in[16:0] >= 8662 && in <= 8671) out = 3654;
	 	 	 else if (in[16:0] >= 8672 && in <= 8681) out = 3655;
	 	 	 else if (in[16:0] >= 8682 && in <= 8692) out = 3656;
	 	 	 else if (in[16:0] >= 8693 && in <= 8702) out = 3657;
	 	 	 else if (in[16:0] >= 8703 && in <= 8713) out = 3658;
	 	 	 else if (in[16:0] >= 8714 && in <= 8723) out = 3659;
	 	 	 else if (in[16:0] >= 8724 && in <= 8734) out = 3660;
	 	 	 else if (in[16:0] >= 8735 && in <= 8745) out = 3661;
	 	 	 else if (in[16:0] >= 8746 && in <= 8755) out = 3662;
	 	 	 else if (in[16:0] >= 8756 && in <= 8766) out = 3663;
	 	 	 else if (in[16:0] >= 8767 && in <= 8776) out = 3664;
	 	 	 else if (in[16:0] >= 8777 && in <= 8787) out = 3665;
	 	 	 else if (in[16:0] >= 8788 && in <= 8798) out = 3666;
	 	 	 else if (in[16:0] >= 8799 && in <= 8808) out = 3667;
	 	 	 else if (in[16:0] >= 8809 && in <= 8819) out = 3668;
	 	 	 else if (in[16:0] >= 8820 && in <= 8830) out = 3669;
	 	 	 else if (in[16:0] >= 8831 && in <= 8841) out = 3670;
	 	 	 else if (in[16:0] >= 8842 && in <= 8851) out = 3671;
	 	 	 else if (in[16:0] >= 8852 && in <= 8862) out = 3672;
	 	 	 else if (in[16:0] >= 8863 && in <= 8873) out = 3673;
	 	 	 else if (in[16:0] >= 8874 && in <= 8884) out = 3674;
	 	 	 else if (in[16:0] >= 8885 && in <= 8895) out = 3675;
	 	 	 else if (in[16:0] >= 8896 && in <= 8906) out = 3676;
	 	 	 else if (in[16:0] >= 8907 && in <= 8917) out = 3677;
	 	 	 else if (in[16:0] >= 8918 && in <= 8928) out = 3678;
	 	 	 else if (in[16:0] >= 8929 && in <= 8939) out = 3679;
	 	 	 else if (in[16:0] >= 8940 && in <= 8950) out = 3680;
	 	 	 else if (in[16:0] >= 8951 && in <= 8961) out = 3681;
	 	 	 else if (in[16:0] >= 8962 && in <= 8972) out = 3682;
	 	 	 else if (in[16:0] >= 8973 && in <= 8983) out = 3683;
	 	 	 else if (in[16:0] >= 8984 && in <= 8994) out = 3684;
	 	 	 else if (in[16:0] >= 8995 && in <= 9005) out = 3685;
	 	 	 else if (in[16:0] >= 9006 && in <= 9016) out = 3686;
	 	 	 else if (in[16:0] >= 9017 && in <= 9027) out = 3687;
	 	 	 else if (in[16:0] >= 9028 && in <= 9038) out = 3688;
	 	 	 else if (in[16:0] >= 9039 && in <= 9050) out = 3689;
	 	 	 else if (in[16:0] >= 9051 && in <= 9061) out = 3690;
	 	 	 else if (in[16:0] >= 9062 && in <= 9072) out = 3691;
	 	 	 else if (in[16:0] >= 9073 && in <= 9083) out = 3692;
	 	 	 else if (in[16:0] >= 9084 && in <= 9095) out = 3693;
	 	 	 else if (in[16:0] >= 9096 && in <= 9106) out = 3694;
	 	 	 else if (in[16:0] >= 9107 && in <= 9117) out = 3695;
	 	 	 else if (in[16:0] >= 9118 && in <= 9129) out = 3696;
	 	 	 else if (in[16:0] >= 9130 && in <= 9140) out = 3697;
	 	 	 else if (in[16:0] >= 9141 && in <= 9152) out = 3698;
	 	 	 else if (in[16:0] >= 9153 && in <= 9163) out = 3699;
	 	 	 else if (in[16:0] >= 9164 && in <= 9175) out = 3700;
	 	 	 else if (in[16:0] >= 9176 && in <= 9186) out = 3701;
	 	 	 else if (in[16:0] >= 9187 && in <= 9198) out = 3702;
	 	 	 else if (in[16:0] >= 9199 && in <= 9209) out = 3703;
	 	 	 else if (in[16:0] >= 9210 && in <= 9221) out = 3704;
	 	 	 else if (in[16:0] >= 9222 && in <= 9232) out = 3705;
	 	 	 else if (in[16:0] >= 9233 && in <= 9244) out = 3706;
	 	 	 else if (in[16:0] >= 9245 && in <= 9256) out = 3707;
	 	 	 else if (in[16:0] >= 9257 && in <= 9267) out = 3708;
	 	 	 else if (in[16:0] >= 9268 && in <= 9279) out = 3709;
	 	 	 else if (in[16:0] >= 9280 && in <= 9291) out = 3710;
	 	 	 else if (in[16:0] >= 9292 && in <= 9303) out = 3711;
	 	 	 else if (in[16:0] >= 9304 && in <= 9315) out = 3712;
	 	 	 else if (in[16:0] >= 9316 && in <= 9326) out = 3713;
	 	 	 else if (in[16:0] >= 9327 && in <= 9338) out = 3714;
	 	 	 else if (in[16:0] >= 9339 && in <= 9350) out = 3715;
	 	 	 else if (in[16:0] >= 9351 && in <= 9362) out = 3716;
	 	 	 else if (in[16:0] >= 9363 && in <= 9374) out = 3717;
	 	 	 else if (in[16:0] >= 9375 && in <= 9386) out = 3718;
	 	 	 else if (in[16:0] >= 9387 && in <= 9398) out = 3719;
	 	 	 else if (in[16:0] >= 9399 && in <= 9410) out = 3720;
	 	 	 else if (in[16:0] >= 9411 && in <= 9422) out = 3721;
	 	 	 else if (in[16:0] >= 9423 && in <= 9434) out = 3722;
	 	 	 else if (in[16:0] >= 9435 && in <= 9446) out = 3723;
	 	 	 else if (in[16:0] >= 9447 && in <= 9458) out = 3724;
	 	 	 else if (in[16:0] >= 9459 && in <= 9471) out = 3725;
	 	 	 else if (in[16:0] >= 9472 && in <= 9483) out = 3726;
	 	 	 else if (in[16:0] >= 9484 && in <= 9495) out = 3727;
	 	 	 else if (in[16:0] >= 9496 && in <= 9507) out = 3728;
	 	 	 else if (in[16:0] >= 9508 && in <= 9520) out = 3729;
	 	 	 else if (in[16:0] >= 9521 && in <= 9532) out = 3730;
	 	 	 else if (in[16:0] >= 9533 && in <= 9544) out = 3731;
	 	 	 else if (in[16:0] >= 9545 && in <= 9557) out = 3732;
	 	 	 else if (in[16:0] >= 9558 && in <= 9569) out = 3733;
	 	 	 else if (in[16:0] >= 9570 && in <= 9582) out = 3734;
	 	 	 else if (in[16:0] >= 9583 && in <= 9594) out = 3735;
	 	 	 else if (in[16:0] >= 9595 && in <= 9607) out = 3736;
	 	 	 else if (in[16:0] >= 9608 && in <= 9619) out = 3737;
	 	 	 else if (in[16:0] >= 9620 && in <= 9632) out = 3738;
	 	 	 else if (in[16:0] >= 9633 && in <= 9644) out = 3739;
	 	 	 else if (in[16:0] >= 9645 && in <= 9657) out = 3740;
	 	 	 else if (in[16:0] >= 9658 && in <= 9670) out = 3741;
	 	 	 else if (in[16:0] >= 9671 && in <= 9682) out = 3742;
	 	 	 else if (in[16:0] >= 9683 && in <= 9695) out = 3743;
	 	 	 else if (in[16:0] >= 9696 && in <= 9708) out = 3744;
	 	 	 else if (in[16:0] >= 9709 && in <= 9721) out = 3745;
	 	 	 else if (in[16:0] >= 9722 && in <= 9734) out = 3746;
	 	 	 else if (in[16:0] >= 9735 && in <= 9747) out = 3747;
	 	 	 else if (in[16:0] >= 9748 && in <= 9759) out = 3748;
	 	 	 else if (in[16:0] >= 9760 && in <= 9772) out = 3749;
	 	 	 else if (in[16:0] >= 9773 && in <= 9785) out = 3750;
	 	 	 else if (in[16:0] >= 9786 && in <= 9798) out = 3751;
	 	 	 else if (in[16:0] >= 9799 && in <= 9811) out = 3752;
	 	 	 else if (in[16:0] >= 9812 && in <= 9825) out = 3753;
	 	 	 else if (in[16:0] >= 9826 && in <= 9838) out = 3754;
	 	 	 else if (in[16:0] >= 9839 && in <= 9851) out = 3755;
	 	 	 else if (in[16:0] >= 9852 && in <= 9864) out = 3756;
	 	 	 else if (in[16:0] >= 9865 && in <= 9877) out = 3757;
	 	 	 else if (in[16:0] >= 9878 && in <= 9891) out = 3758;
	 	 	 else if (in[16:0] >= 9892 && in <= 9904) out = 3759;
	 	 	 else if (in[16:0] >= 9905 && in <= 9917) out = 3760;
	 	 	 else if (in[16:0] >= 9918 && in <= 9931) out = 3761;
	 	 	 else if (in[16:0] >= 9932 && in <= 9944) out = 3762;
	 	 	 else if (in[16:0] >= 9945 && in <= 9957) out = 3763;
	 	 	 else if (in[16:0] >= 9958 && in <= 9971) out = 3764;
	 	 	 else if (in[16:0] >= 9972 && in <= 9984) out = 3765;
	 	 	 else if (in[16:0] >= 9985 && in <= 9998) out = 3766;
	 	 	 else if (in[16:0] >= 9999 && in <= 10012) out = 3767;
	 	 	 else if (in[16:0] >= 10013 && in <= 10025) out = 3768;
	 	 	 else if (in[16:0] >= 10026 && in <= 10039) out = 3769;
	 	 	 else if (in[16:0] >= 10040 && in <= 10053) out = 3770;
	 	 	 else if (in[16:0] >= 10054 && in <= 10066) out = 3771;
	 	 	 else if (in[16:0] >= 10067 && in <= 10080) out = 3772;
	 	 	 else if (in[16:0] >= 10081 && in <= 10094) out = 3773;
	 	 	 else if (in[16:0] >= 10095 && in <= 10108) out = 3774;
	 	 	 else if (in[16:0] >= 10109 && in <= 10122) out = 3775;
	 	 	 else if (in[16:0] >= 10123 && in <= 10136) out = 3776;
	 	 	 else if (in[16:0] >= 10137 && in <= 10150) out = 3777;
	 	 	 else if (in[16:0] >= 10151 && in <= 10164) out = 3778;
	 	 	 else if (in[16:0] >= 10165 && in <= 10178) out = 3779;
	 	 	 else if (in[16:0] >= 10179 && in <= 10192) out = 3780;
	 	 	 else if (in[16:0] >= 10193 && in <= 10206) out = 3781;
	 	 	 else if (in[16:0] >= 10207 && in <= 10220) out = 3782;
	 	 	 else if (in[16:0] >= 10221 && in <= 10234) out = 3783;
	 	 	 else if (in[16:0] >= 10235 && in <= 10249) out = 3784;
	 	 	 else if (in[16:0] >= 10250 && in <= 10263) out = 3785;
	 	 	 else if (in[16:0] >= 10264 && in <= 10277) out = 3786;
	 	 	 else if (in[16:0] >= 10278 && in <= 10292) out = 3787;
	 	 	 else if (in[16:0] >= 10293 && in <= 10306) out = 3788;
	 	 	 else if (in[16:0] >= 10307 && in <= 10321) out = 3789;
	 	 	 else if (in[16:0] >= 10322 && in <= 10335) out = 3790;
	 	 	 else if (in[16:0] >= 10336 && in <= 10350) out = 3791;
	 	 	 else if (in[16:0] >= 10351 && in <= 10364) out = 3792;
	 	 	 else if (in[16:0] >= 10365 && in <= 10379) out = 3793;
	 	 	 else if (in[16:0] >= 10380 && in <= 10394) out = 3794;
	 	 	 else if (in[16:0] >= 10395 && in <= 10408) out = 3795;
	 	 	 else if (in[16:0] >= 10409 && in <= 10423) out = 3796;
	 	 	 else if (in[16:0] >= 10424 && in <= 10438) out = 3797;
	 	 	 else if (in[16:0] >= 10439 && in <= 10453) out = 3798;
	 	 	 else if (in[16:0] >= 10454 && in <= 10468) out = 3799;
	 	 	 else if (in[16:0] >= 10469 && in <= 10483) out = 3800;
	 	 	 else if (in[16:0] >= 10484 && in <= 10498) out = 3801;
	 	 	 else if (in[16:0] >= 10499 && in <= 10513) out = 3802;
	 	 	 else if (in[16:0] >= 10514 && in <= 10528) out = 3803;
	 	 	 else if (in[16:0] >= 10529 && in <= 10543) out = 3804;
	 	 	 else if (in[16:0] >= 10544 && in <= 10559) out = 3805;
	 	 	 else if (in[16:0] >= 10560 && in <= 10574) out = 3806;
	 	 	 else if (in[16:0] >= 10575 && in <= 10589) out = 3807;
	 	 	 else if (in[16:0] >= 10590 && in <= 10605) out = 3808;
	 	 	 else if (in[16:0] >= 10606 && in <= 10620) out = 3809;
	 	 	 else if (in[16:0] >= 10621 && in <= 10635) out = 3810;
	 	 	 else if (in[16:0] >= 10636 && in <= 10651) out = 3811;
	 	 	 else if (in[16:0] >= 10652 && in <= 10667) out = 3812;
	 	 	 else if (in[16:0] >= 10668 && in <= 10682) out = 3813;
	 	 	 else if (in[16:0] >= 10683 && in <= 10698) out = 3814;
	 	 	 else if (in[16:0] >= 10699 && in <= 10714) out = 3815;
	 	 	 else if (in[16:0] >= 10715 && in <= 10729) out = 3816;
	 	 	 else if (in[16:0] >= 10730 && in <= 10745) out = 3817;
	 	 	 else if (in[16:0] >= 10746 && in <= 10761) out = 3818;
	 	 	 else if (in[16:0] >= 10762 && in <= 10777) out = 3819;
	 	 	 else if (in[16:0] >= 10778 && in <= 10793) out = 3820;
	 	 	 else if (in[16:0] >= 10794 && in <= 10809) out = 3821;
	 	 	 else if (in[16:0] >= 10810 && in <= 10825) out = 3822;
	 	 	 else if (in[16:0] >= 10826 && in <= 10841) out = 3823;
	 	 	 else if (in[16:0] >= 10842 && in <= 10858) out = 3824;
	 	 	 else if (in[16:0] >= 10859 && in <= 10874) out = 3825;
	 	 	 else if (in[16:0] >= 10875 && in <= 10890) out = 3826;
	 	 	 else if (in[16:0] >= 10891 && in <= 10907) out = 3827;
	 	 	 else if (in[16:0] >= 10908 && in <= 10923) out = 3828;
	 	 	 else if (in[16:0] >= 10924 && in <= 10939) out = 3829;
	 	 	 else if (in[16:0] >= 10940 && in <= 10956) out = 3830;
	 	 	 else if (in[16:0] >= 10957 && in <= 10973) out = 3831;
	 	 	 else if (in[16:0] >= 10974 && in <= 10989) out = 3832;
	 	 	 else if (in[16:0] >= 10990 && in <= 11006) out = 3833;
	 	 	 else if (in[16:0] >= 11007 && in <= 11023) out = 3834;
	 	 	 else if (in[16:0] >= 11024 && in <= 11040) out = 3835;
	 	 	 else if (in[16:0] >= 11041 && in <= 11057) out = 3836;
	 	 	 else if (in[16:0] >= 11058 && in <= 11074) out = 3837;
	 	 	 else if (in[16:0] >= 11075 && in <= 11091) out = 3838;
	 	 	 else if (in[16:0] >= 11092 && in <= 11108) out = 3839;
	 	 	 else if (in[16:0] >= 11109 && in <= 11125) out = 3840;
	 	 	 else if (in[16:0] >= 11126 && in <= 11142) out = 3841;
	 	 	 else if (in[16:0] >= 11143 && in <= 11159) out = 3842;
	 	 	 else if (in[16:0] >= 11160 && in <= 11177) out = 3843;
	 	 	 else if (in[16:0] >= 11178 && in <= 11194) out = 3844;
	 	 	 else if (in[16:0] >= 11195 && in <= 11212) out = 3845;
	 	 	 else if (in[16:0] >= 11213 && in <= 11229) out = 3846;
	 	 	 else if (in[16:0] >= 11230 && in <= 11247) out = 3847;
	 	 	 else if (in[16:0] >= 11248 && in <= 11264) out = 3848;
	 	 	 else if (in[16:0] >= 11265 && in <= 11282) out = 3849;
	 	 	 else if (in[16:0] >= 11283 && in <= 11300) out = 3850;
	 	 	 else if (in[16:0] >= 11301 && in <= 11318) out = 3851;
	 	 	 else if (in[16:0] >= 11319 && in <= 11336) out = 3852;
	 	 	 else if (in[16:0] >= 11337 && in <= 11354) out = 3853;
	 	 	 else if (in[16:0] >= 11355 && in <= 11372) out = 3854;
	 	 	 else if (in[16:0] >= 11373 && in <= 11390) out = 3855;
	 	 	 else if (in[16:0] >= 11391 && in <= 11408) out = 3856;
	 	 	 else if (in[16:0] >= 11409 && in <= 11427) out = 3857;
	 	 	 else if (in[16:0] >= 11428 && in <= 11445) out = 3858;
	 	 	 else if (in[16:0] >= 11446 && in <= 11464) out = 3859;
	 	 	 else if (in[16:0] >= 11465 && in <= 11482) out = 3860;
	 	 	 else if (in[16:0] >= 11483 && in <= 11501) out = 3861;
	 	 	 else if (in[16:0] >= 11502 && in <= 11519) out = 3862;
	 	 	 else if (in[16:0] >= 11520 && in <= 11538) out = 3863;
	 	 	 else if (in[16:0] >= 11539 && in <= 11557) out = 3864;
	 	 	 else if (in[16:0] >= 11558 && in <= 11576) out = 3865;
	 	 	 else if (in[16:0] >= 11577 && in <= 11595) out = 3866;
	 	 	 else if (in[16:0] >= 11596 && in <= 11614) out = 3867;
	 	 	 else if (in[16:0] >= 11615 && in <= 11633) out = 3868;
	 	 	 else if (in[16:0] >= 11634 && in <= 11652) out = 3869;
	 	 	 else if (in[16:0] >= 11653 && in <= 11672) out = 3870;
	 	 	 else if (in[16:0] >= 11673 && in <= 11691) out = 3871;
	 	 	 else if (in[16:0] >= 11692 && in <= 11710) out = 3872;
	 	 	 else if (in[16:0] >= 11711 && in <= 11730) out = 3873;
	 	 	 else if (in[16:0] >= 11731 && in <= 11750) out = 3874;
	 	 	 else if (in[16:0] >= 11751 && in <= 11769) out = 3875;
	 	 	 else if (in[16:0] >= 11770 && in <= 11789) out = 3876;
	 	 	 else if (in[16:0] >= 11790 && in <= 11809) out = 3877;
	 	 	 else if (in[16:0] >= 11810 && in <= 11829) out = 3878;
	 	 	 else if (in[16:0] >= 11830 && in <= 11849) out = 3879;
	 	 	 else if (in[16:0] >= 11850 && in <= 11869) out = 3880;
	 	 	 else if (in[16:0] >= 11870 && in <= 11889) out = 3881;
	 	 	 else if (in[16:0] >= 11890 && in <= 11910) out = 3882;
	 	 	 else if (in[16:0] >= 11911 && in <= 11930) out = 3883;
	 	 	 else if (in[16:0] >= 11931 && in <= 11951) out = 3884;
	 	 	 else if (in[16:0] >= 11952 && in <= 11971) out = 3885;
	 	 	 else if (in[16:0] >= 11972 && in <= 11992) out = 3886;
	 	 	 else if (in[16:0] >= 11993 && in <= 12013) out = 3887;
	 	 	 else if (in[16:0] >= 12014 && in <= 12034) out = 3888;
	 	 	 else if (in[16:0] >= 12035 && in <= 12055) out = 3889;
	 	 	 else if (in[16:0] >= 12056 && in <= 12076) out = 3890;
	 	 	 else if (in[16:0] >= 12077 && in <= 12097) out = 3891;
	 	 	 else if (in[16:0] >= 12098 && in <= 12118) out = 3892;
	 	 	 else if (in[16:0] >= 12119 && in <= 12140) out = 3893;
	 	 	 else if (in[16:0] >= 12141 && in <= 12161) out = 3894;
	 	 	 else if (in[16:0] >= 12162 && in <= 12183) out = 3895;
	 	 	 else if (in[16:0] >= 12184 && in <= 12204) out = 3896;
	 	 	 else if (in[16:0] >= 12205 && in <= 12226) out = 3897;
	 	 	 else if (in[16:0] >= 12227 && in <= 12248) out = 3898;
	 	 	 else if (in[16:0] >= 12249 && in <= 12270) out = 3899;
	 	 	 else if (in[16:0] >= 12271 && in <= 12292) out = 3900;
	 	 	 else if (in[16:0] >= 12293 && in <= 12314) out = 3901;
	 	 	 else if (in[16:0] >= 12315 && in <= 12337) out = 3902;
	 	 	 else if (in[16:0] >= 12338 && in <= 12359) out = 3903;
	 	 	 else if (in[16:0] >= 12360 && in <= 12382) out = 3904;
	 	 	 else if (in[16:0] >= 12383 && in <= 12404) out = 3905;
	 	 	 else if (in[16:0] >= 12405 && in <= 12427) out = 3906;
	 	 	 else if (in[16:0] >= 12428 && in <= 12450) out = 3907;
	 	 	 else if (in[16:0] >= 12451 && in <= 12473) out = 3908;
	 	 	 else if (in[16:0] >= 12474 && in <= 12496) out = 3909;
	 	 	 else if (in[16:0] >= 12497 && in <= 12519) out = 3910;
	 	 	 else if (in[16:0] >= 12520 && in <= 12543) out = 3911;
	 	 	 else if (in[16:0] >= 12544 && in <= 12566) out = 3912;
	 	 	 else if (in[16:0] >= 12567 && in <= 12590) out = 3913;
	 	 	 else if (in[16:0] >= 12591 && in <= 12614) out = 3914;
	 	 	 else if (in[16:0] >= 12615 && in <= 12637) out = 3915;
	 	 	 else if (in[16:0] >= 12638 && in <= 12661) out = 3916;
	 	 	 else if (in[16:0] >= 12662 && in <= 12686) out = 3917;
	 	 	 else if (in[16:0] >= 12687 && in <= 12710) out = 3918;
	 	 	 else if (in[16:0] >= 12711 && in <= 12734) out = 3919;
	 	 	 else if (in[16:0] >= 12735 && in <= 12759) out = 3920;
	 	 	 else if (in[16:0] >= 12760 && in <= 12783) out = 3921;
	 	 	 else if (in[16:0] >= 12784 && in <= 12808) out = 3922;
	 	 	 else if (in[16:0] >= 12809 && in <= 12833) out = 3923;
	 	 	 else if (in[16:0] >= 12834 && in <= 12858) out = 3924;
	 	 	 else if (in[16:0] >= 12859 && in <= 12883) out = 3925;
	 	 	 else if (in[16:0] >= 12884 && in <= 12909) out = 3926;
	 	 	 else if (in[16:0] >= 12910 && in <= 12934) out = 3927;
	 	 	 else if (in[16:0] >= 12935 && in <= 12960) out = 3928;
	 	 	 else if (in[16:0] >= 12961 && in <= 12986) out = 3929;
	 	 	 else if (in[16:0] >= 12987 && in <= 13012) out = 3930;
	 	 	 else if (in[16:0] >= 13013 && in <= 13038) out = 3931;
	 	 	 else if (in[16:0] >= 13039 && in <= 13064) out = 3932;
	 	 	 else if (in[16:0] >= 13065 && in <= 13090) out = 3933;
	 	 	 else if (in[16:0] >= 13091 && in <= 13117) out = 3934;
	 	 	 else if (in[16:0] >= 13118 && in <= 13144) out = 3935;
	 	 	 else if (in[16:0] >= 13145 && in <= 13171) out = 3936;
	 	 	 else if (in[16:0] >= 13172 && in <= 13198) out = 3937;
	 	 	 else if (in[16:0] >= 13199 && in <= 13225) out = 3938;
	 	 	 else if (in[16:0] >= 13226 && in <= 13252) out = 3939;
	 	 	 else if (in[16:0] >= 13253 && in <= 13280) out = 3940;
	 	 	 else if (in[16:0] >= 13281 && in <= 13307) out = 3941;
	 	 	 else if (in[16:0] >= 13308 && in <= 13335) out = 3942;
	 	 	 else if (in[16:0] >= 13336 && in <= 13363) out = 3943;
	 	 	 else if (in[16:0] >= 13364 && in <= 13392) out = 3944;
	 	 	 else if (in[16:0] >= 13393 && in <= 13420) out = 3945;
	 	 	 else if (in[16:0] >= 13421 && in <= 13449) out = 3946;
	 	 	 else if (in[16:0] >= 13450 && in <= 13478) out = 3947;
	 	 	 else if (in[16:0] >= 13479 && in <= 13507) out = 3948;
	 	 	 else if (in[16:0] >= 13508 && in <= 13536) out = 3949;
	 	 	 else if (in[16:0] >= 13537 && in <= 13565) out = 3950;
	 	 	 else if (in[16:0] >= 13566 && in <= 13595) out = 3951;
	 	 	 else if (in[16:0] >= 13596 && in <= 13624) out = 3952;
	 	 	 else if (in[16:0] >= 13625 && in <= 13654) out = 3953;
	 	 	 else if (in[16:0] >= 13655 && in <= 13685) out = 3954;
	 	 	 else if (in[16:0] >= 13686 && in <= 13715) out = 3955;
	 	 	 else if (in[16:0] >= 13716 && in <= 13746) out = 3956;
	 	 	 else if (in[16:0] >= 13747 && in <= 13776) out = 3957;
	 	 	 else if (in[16:0] >= 13777 && in <= 13807) out = 3958;
	 	 	 else if (in[16:0] >= 13808 && in <= 13839) out = 3959;
	 	 	 else if (in[16:0] >= 13840 && in <= 13870) out = 3960;
	 	 	 else if (in[16:0] >= 13871 && in <= 13902) out = 3961;
	 	 	 else if (in[16:0] >= 13903 && in <= 13934) out = 3962;
	 	 	 else if (in[16:0] >= 13935 && in <= 13966) out = 3963;
	 	 	 else if (in[16:0] >= 13967 && in <= 13999) out = 3964;
	 	 	 else if (in[16:0] >= 14000 && in <= 14031) out = 3965;
	 	 	 else if (in[16:0] >= 14032 && in <= 14064) out = 3966;
	 	 	 else if (in[16:0] >= 14065 && in <= 14097) out = 3967;
	 	 	 else if (in[16:0] >= 14098 && in <= 14131) out = 3968;
	 	 	 else if (in[16:0] >= 14132 && in <= 14164) out = 3969;
	 	 	 else if (in[16:0] >= 14165 && in <= 14198) out = 3970;
	 	 	 else if (in[16:0] >= 14199 && in <= 14232) out = 3971;
	 	 	 else if (in[16:0] >= 14233 && in <= 14267) out = 3972;
	 	 	 else if (in[16:0] >= 14268 && in <= 14302) out = 3973;
	 	 	 else if (in[16:0] >= 14303 && in <= 14337) out = 3974;
	 	 	 else if (in[16:0] >= 14338 && in <= 14372) out = 3975;
	 	 	 else if (in[16:0] >= 14373 && in <= 14408) out = 3976;
	 	 	 else if (in[16:0] >= 14409 && in <= 14443) out = 3977;
	 	 	 else if (in[16:0] >= 14444 && in <= 14480) out = 3978;
	 	 	 else if (in[16:0] >= 14481 && in <= 14516) out = 3979;
	 	 	 else if (in[16:0] >= 14517 && in <= 14553) out = 3980;
	 	 	 else if (in[16:0] >= 14554 && in <= 14590) out = 3981;
	 	 	 else if (in[16:0] >= 14591 && in <= 14628) out = 3982;
	 	 	 else if (in[16:0] >= 14629 && in <= 14665) out = 3983;
	 	 	 else if (in[16:0] >= 14666 && in <= 14703) out = 3984;
	 	 	 else if (in[16:0] >= 14704 && in <= 14742) out = 3985;
	 	 	 else if (in[16:0] >= 14743 && in <= 14781) out = 3986;
	 	 	 else if (in[16:0] >= 14782 && in <= 14820) out = 3987;
	 	 	 else if (in[16:0] >= 14821 && in <= 14859) out = 3988;
	 	 	 else if (in[16:0] >= 14860 && in <= 14899) out = 3989;
	 	 	 else if (in[16:0] >= 14900 && in <= 14939) out = 3990;
	 	 	 else if (in[16:0] >= 14940 && in <= 14980) out = 3991;
	 	 	 else if (in[16:0] >= 14981 && in <= 15021) out = 3992;
	 	 	 else if (in[16:0] >= 15022 && in <= 15062) out = 3993;
	 	 	 else if (in[16:0] >= 15063 && in <= 15104) out = 3994;
	 	 	 else if (in[16:0] >= 15105 && in <= 15146) out = 3995;
	 	 	 else if (in[16:0] >= 15147 && in <= 15189) out = 3996;
	 	 	 else if (in[16:0] >= 15190 && in <= 15232) out = 3997;
	 	 	 else if (in[16:0] >= 15233 && in <= 15275) out = 3998;
	 	 	 else if (in[16:0] >= 15276 && in <= 15319) out = 3999;
	 	 	 else if (in[16:0] >= 15320 && in <= 15364) out = 4000;
	 	 	 else if (in[16:0] >= 15365 && in <= 15408) out = 4001;
	 	 	 else if (in[16:0] >= 15409 && in <= 15454) out = 4002;
	 	 	 else if (in[16:0] >= 15455 && in <= 15500) out = 4003;
	 	 	 else if (in[16:0] >= 15501 && in <= 15546) out = 4004;
	 	 	 else if (in[16:0] >= 15547 && in <= 15593) out = 4005;
	 	 	 else if (in[16:0] >= 15594 && in <= 15640) out = 4006;
	 	 	 else if (in[16:0] >= 15641 && in <= 15688) out = 4007;
	 	 	 else if (in[16:0] >= 15689 && in <= 15736) out = 4008;
	 	 	 else if (in[16:0] >= 15737 && in <= 15785) out = 4009;
	 	 	 else if (in[16:0] >= 15786 && in <= 15835) out = 4010;
	 	 	 else if (in[16:0] >= 15836 && in <= 15885) out = 4011;
	 	 	 else if (in[16:0] >= 15886 && in <= 15935) out = 4012;
	 	 	 else if (in[16:0] >= 15936 && in <= 15987) out = 4013;
	 	 	 else if (in[16:0] >= 15988 && in <= 16038) out = 4014;
	 	 	 else if (in[16:0] >= 16039 && in <= 16091) out = 4015;
	 	 	 else if (in[16:0] >= 16092 && in <= 16144) out = 4016;
	 	 	 else if (in[16:0] >= 16145 && in <= 16198) out = 4017;
	 	 	 else if (in[16:0] >= 16199 && in <= 16253) out = 4018;
	 	 	 else if (in[16:0] >= 16254 && in <= 16308) out = 4019;
	 	 	 else if (in[16:0] >= 16309 && in <= 16364) out = 4020;
	 	 	 else if (in[16:0] >= 16365 && in <= 16421) out = 4021;
	 	 	 else if (in[16:0] >= 16422 && in <= 16478) out = 4022;
	 	 	 else if (in[16:0] >= 16479 && in <= 16536) out = 4023;
	 	 	 else if (in[16:0] >= 16537 && in <= 16596) out = 4024;
	 	 	 else if (in[16:0] >= 16597 && in <= 16656) out = 4025;
	 	 	 else if (in[16:0] >= 16657 && in <= 16716) out = 4026;
	 	 	 else if (in[16:0] >= 16717 && in <= 16778) out = 4027;
	 	 	 else if (in[16:0] >= 16779 && in <= 16841) out = 4028;
	 	 	 else if (in[16:0] >= 16842 && in <= 16904) out = 4029;
	 	 	 else if (in[16:0] >= 16905 && in <= 16969) out = 4030;
	 	 	 else if (in[16:0] >= 16970 && in <= 17034) out = 4031;
	 	 	 else if (in[16:0] >= 17035 && in <= 17101) out = 4032;
	 	 	 else if (in[16:0] >= 17102 && in <= 17168) out = 4033;
	 	 	 else if (in[16:0] >= 17169 && in <= 17237) out = 4034;
	 	 	 else if (in[16:0] >= 17238 && in <= 17307) out = 4035;
	 	 	 else if (in[16:0] >= 17308 && in <= 17378) out = 4036;
	 	 	 else if (in[16:0] >= 17379 && in <= 17450) out = 4037;
	 	 	 else if (in[16:0] >= 17451 && in <= 17524) out = 4038;
	 	 	 else if (in[16:0] >= 17525 && in <= 17599) out = 4039;
	 	 	 else if (in[16:0] >= 17600 && in <= 17675) out = 4040;
	 	 	 else if (in[16:0] >= 17676 && in <= 17752) out = 4041;
	 	 	 else if (in[16:0] >= 17753 && in <= 17831) out = 4042;
	 	 	 else if (in[16:0] >= 17832 && in <= 17912) out = 4043;
	 	 	 else if (in[16:0] >= 17913 && in <= 17994) out = 4044;
	 	 	 else if (in[16:0] >= 17995 && in <= 18078) out = 4045;
	 	 	 else if (in[16:0] >= 18079 && in <= 18163) out = 4046;
	 	 	 else if (in[16:0] >= 18164 && in <= 18251) out = 4047;
	 	 	 else if (in[16:0] >= 18252 && in <= 18340) out = 4048;
	 	 	 else if (in[16:0] >= 18341 && in <= 18431) out = 4049;
	 	 	 else if (in[16:0] >= 18432 && in <= 18524) out = 4050;
	 	 	 else if (in[16:0] >= 18525 && in <= 18619) out = 4051;
	 	 	 else if (in[16:0] >= 18620 && in <= 18716) out = 4052;
	 	 	 else if (in[16:0] >= 18717 && in <= 18816) out = 4053;
	 	 	 else if (in[16:0] >= 18817 && in <= 18918) out = 4054;
	 	 	 else if (in[16:0] >= 18919 && in <= 19023) out = 4055;
	 	 	 else if (in[16:0] >= 19024 && in <= 19130) out = 4056;
	 	 	 else if (in[16:0] >= 19131 && in <= 19241) out = 4057;
	 	 	 else if (in[16:0] >= 19242 && in <= 19354) out = 4058;
	 	 	 else if (in[16:0] >= 19355 && in <= 19470) out = 4059;
	 	 	 else if (in[16:0] >= 19471 && in <= 19590) out = 4060;
	 	 	 else if (in[16:0] >= 19591 && in <= 19713) out = 4061;
	 	 	 else if (in[16:0] >= 19714 && in <= 19840) out = 4062;
	 	 	 else if (in[16:0] >= 19841 && in <= 19971) out = 4063;
	 	 	 else if (in[16:0] >= 19972 && in <= 20107) out = 4064;
	 	 	 else if (in[16:0] >= 20108 && in <= 20247) out = 4065;
	 	 	 else if (in[16:0] >= 20248 && in <= 20391) out = 4066;
	 	 	 else if (in[16:0] >= 20392 && in <= 20541) out = 4067;
	 	 	 else if (in[16:0] >= 20542 && in <= 20697) out = 4068;
	 	 	 else if (in[16:0] >= 20698 && in <= 20858) out = 4069;
	 	 	 else if (in[16:0] >= 20859 && in <= 21027) out = 4070;
	 	 	 else if (in[16:0] >= 21028 && in <= 21202) out = 4071;
	 	 	 else if (in[16:0] >= 21203 && in <= 21385) out = 4072;
	 	 	 else if (in[16:0] >= 21386 && in <= 21577) out = 4073;
	 	 	 else if (in[16:0] >= 21578 && in <= 21777) out = 4074;
	 	 	 else if (in[16:0] >= 21778 && in <= 21989) out = 4075;
	 	 	 else if (in[16:0] >= 21990 && in <= 22211) out = 4076;
	 	 	 else if (in[16:0] >= 22212 && in <= 22446) out = 4077;
	 	 	 else if (in[16:0] >= 22447 && in <= 22696) out = 4078;
	 	 	 else if (in[16:0] >= 22697 && in <= 22961) out = 4079;
	 	 	 else if (in[16:0] >= 22962 && in <= 23244) out = 4080;
	 	 	 else if (in[16:0] >= 23245 && in <= 23549) out = 4081;
	 	 	 else if (in[16:0] >= 23550 && in <= 23878) out = 4082;
	 	 	 else if (in[16:0] >= 23879 && in <= 24235) out = 4083;
	 	 	 else if (in[16:0] >= 24236 && in <= 24627) out = 4084;
	 	 	 else if (in[16:0] >= 24628 && in <= 25059) out = 4085;
	 	 	 else if (in[16:0] >= 25060 && in <= 25543) out = 4086;
	 	 	 else if (in[16:0] >= 25544 && in <= 26091) out = 4087;
	 	 	 else if (in[16:0] >= 26092 && in <= 26723) out = 4088;
	 	 	 else if (in[16:0] >= 26724 && in <= 27471) out = 4089;
	 	 	 else if (in[16:0] >= 27472 && in <= 28386) out = 4090;
	 	 	 else if (in[16:0] >= 28387 && in <= 29565) out = 4091;
	 	 	 else if (in[16:0] >= 29566 && in <= 31227) out = 4092;
	 	 	 else if (in[16:0] >= 31228 && in <= 34067) out = 4093;
	 	 	 else if (in[16:0] >= 34068 && in <= 65535) out = 4094;
	 	 	else out=4095;
	 endmodule
	 */

module sigma_int(input data_type in,
    input logic clk,
	 output data_type out);
	 
	 BRAM_wrapper BRAM_sigma_int(.addra_0(in[15:0]), .clka_0(clk), .douta_0(out[11:0]));
	 
	 assign out[31:12] = 0;
	 
endmodule	 
	 
