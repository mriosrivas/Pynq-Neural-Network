`ifndef typedef
`define typedef
    typedef logic signed [31:0] data_type;
    typedef logic signed [31:0] double_data_type;
`endif

