`include "typedef.vh"


module cross_entropy_table_2(input data_type in,
	 output data_type out);
	 	 always_comb
	 	 	 if (in >= 0 && in <= 1) out = -4096;
	 	 	 else if (in >= 2 && in <= 2) out = -2048;
	 	 	 else if (in >= 3 && in <= 3) out = -1365;
	 	 	 else if (in >= 4 && in <= 4) out = -1024;
	 	 	 else if (in >= 5 && in <= 5) out = -819;
	 	 	 else if (in >= 6 && in <= 6) out = -682;
	 	 	 else if (in >= 7 && in <= 7) out = -585;
	 	 	 else if (in >= 8 && in <= 8) out = -512;
	 	 	 else if (in >= 9 && in <= 9) out = -455;
	 	 	 else if (in >= 10 && in <= 10) out = -409;
	 	 	 else if (in >= 11 && in <= 11) out = -372;
	 	 	 else if (in >= 12 && in <= 12) out = -341;
	 	 	 else if (in >= 13 && in <= 13) out = -315;
	 	 	 else if (in >= 14 && in <= 14) out = -292;
	 	 	 else if (in >= 15 && in <= 15) out = -273;
	 	 	 else if (in >= 16 && in <= 16) out = -256;
	 	 	 else if (in >= 17 && in <= 17) out = -240;
	 	 	 else if (in >= 18 && in <= 18) out = -227;
	 	 	 else if (in >= 19 && in <= 19) out = -215;
	 	 	 else if (in >= 20 && in <= 20) out = -204;
	 	 	 else if (in >= 21 && in <= 21) out = -195;
	 	 	 else if (in >= 22 && in <= 22) out = -186;
	 	 	 else if (in >= 23 && in <= 23) out = -178;
	 	 	 else if (in >= 24 && in <= 24) out = -170;
	 	 	 else if (in >= 25 && in <= 25) out = -163;
	 	 	 else if (in >= 26 && in <= 26) out = -157;
	 	 	 else if (in >= 27 && in <= 27) out = -151;
	 	 	 else if (in >= 28 && in <= 28) out = -146;
	 	 	 else if (in >= 29 && in <= 29) out = -141;
	 	 	 else if (in >= 30 && in <= 30) out = -136;
	 	 	 else if (in >= 31 && in <= 31) out = -132;
	 	 	 else if (in >= 32 && in <= 32) out = -128;
	 	 	 else if (in >= 33 && in <= 33) out = -124;
	 	 	 else if (in >= 34 && in <= 34) out = -120;
	 	 	 else if (in >= 35 && in <= 35) out = -117;
	 	 	 else if (in >= 36 && in <= 36) out = -113;
	 	 	 else if (in >= 37 && in <= 37) out = -110;
	 	 	 else if (in >= 38 && in <= 38) out = -107;
	 	 	 else if (in >= 39 && in <= 39) out = -105;
	 	 	 else if (in >= 40 && in <= 40) out = -102;
	 	 	 else if (in >= 41 && in <= 41) out = -99;
	 	 	 else if (in >= 42 && in <= 42) out = -97;
	 	 	 else if (in >= 43 && in <= 43) out = -95;
	 	 	 else if (in >= 44 && in <= 44) out = -93;
	 	 	 else if (in >= 45 && in <= 45) out = -91;
	 	 	 else if (in >= 46 && in <= 46) out = -89;
	 	 	 else if (in >= 47 && in <= 47) out = -87;
	 	 	 else if (in >= 48 && in <= 48) out = -85;
	 	 	 else if (in >= 49 && in <= 49) out = -83;
	 	 	 else if (in >= 50 && in <= 50) out = -81;
	 	 	 else if (in >= 51 && in <= 51) out = -80;
	 	 	 else if (in >= 52 && in <= 52) out = -78;
	 	 	 else if (in >= 53 && in <= 53) out = -77;
	 	 	 else if (in >= 54 && in <= 54) out = -75;
	 	 	 else if (in >= 55 && in <= 55) out = -74;
	 	 	 else if (in >= 56 && in <= 56) out = -73;
	 	 	 else if (in >= 57 && in <= 57) out = -71;
	 	 	 else if (in >= 58 && in <= 58) out = -70;
	 	 	 else if (in >= 59 && in <= 59) out = -69;
	 	 	 else if (in >= 60 && in <= 60) out = -68;
	 	 	 else if (in >= 61 && in <= 61) out = -67;
	 	 	 else if (in >= 62 && in <= 62) out = -66;
	 	 	 else if (in >= 63 && in <= 63) out = -65;
	 	 	 else if (in >= 64 && in <= 64) out = -64;
	 	 	 else if (in >= 65 && in <= 65) out = -63;
	 	 	 else if (in >= 66 && in <= 66) out = -62;
	 	 	 else if (in >= 67 && in <= 67) out = -61;
	 	 	 else if (in >= 68 && in <= 68) out = -60;
	 	 	 else if (in >= 69 && in <= 69) out = -59;
	 	 	 else if (in >= 70 && in <= 70) out = -58;
	 	 	 else if (in >= 71 && in <= 71) out = -57;
	 	 	 else if (in >= 72 && in <= 73) out = -56;
	 	 	 else if (in >= 74 && in <= 74) out = -55;
	 	 	 else if (in >= 75 && in <= 75) out = -54;
	 	 	 else if (in >= 76 && in <= 77) out = -53;
	 	 	 else if (in >= 78 && in <= 78) out = -52;
	 	 	 else if (in >= 79 && in <= 80) out = -51;
	 	 	 else if (in >= 81 && in <= 81) out = -50;
	 	 	 else if (in >= 82 && in <= 83) out = -49;
	 	 	 else if (in >= 84 && in <= 85) out = -48;
	 	 	 else if (in >= 86 && in <= 87) out = -47;
	 	 	 else if (in >= 88 && in <= 89) out = -46;
	 	 	 else if (in >= 90 && in <= 91) out = -45;
	 	 	 else if (in >= 92 && in <= 93) out = -44;
	 	 	 else if (in >= 94 && in <= 95) out = -43;
	 	 	 else if (in >= 96 && in <= 97) out = -42;
	 	 	 else if (in >= 98 && in <= 99) out = -41;
	 	 	 else if (in >= 100 && in <= 102) out = -40;
	 	 	 else if (in >= 103 && in <= 105) out = -39;
	 	 	 else if (in >= 106 && in <= 107) out = -38;
	 	 	 else if (in >= 108 && in <= 110) out = -37;
	 	 	 else if (in >= 111 && in <= 113) out = -36;
	 	 	 else if (in >= 114 && in <= 117) out = -35;
	 	 	 else if (in >= 118 && in <= 120) out = -34;
	 	 	 else if (in >= 121 && in <= 124) out = -33;
	 	 	 else if (in >= 125 && in <= 128) out = -32;
	 	 	 else if (in >= 129 && in <= 132) out = -31;
	 	 	 else if (in >= 133 && in <= 136) out = -30;
	 	 	 else if (in >= 137 && in <= 141) out = -29;
	 	 	 else if (in >= 142 && in <= 146) out = -28;
	 	 	 else if (in >= 147 && in <= 151) out = -27;
	 	 	 else if (in >= 152 && in <= 157) out = -26;
	 	 	 else if (in >= 158 && in <= 163) out = -25;
	 	 	 else if (in >= 164 && in <= 170) out = -24;
	 	 	 else if (in >= 171 && in <= 178) out = -23;
	 	 	 else if (in >= 179 && in <= 186) out = -22;
	 	 	 else if (in >= 187 && in <= 195) out = -21;
	 	 	 else if (in >= 196 && in <= 204) out = -20;
	 	 	 else if (in >= 205 && in <= 215) out = -19;
	 	 	 else if (in >= 216 && in <= 227) out = -18;
	 	 	 else if (in >= 228 && in <= 240) out = -17;
	 	 	 else if (in >= 241 && in <= 256) out = -16;
	 	 	 else if (in >= 257 && in <= 273) out = -15;
	 	 	 else if (in >= 274 && in <= 292) out = -14;
	 	 	 else if (in >= 293 && in <= 315) out = -13;
	 	 	 else if (in >= 316 && in <= 341) out = -12;
	 	 	 else if (in >= 342 && in <= 372) out = -11;
	 	 	 else if (in >= 373 && in <= 409) out = -10;
	 	 	 else if (in >= 410 && in <= 455) out = -9;
	 	 	 else if (in >= 456 && in <= 512) out = -8;
	 	 	 else if (in >= 513 && in <= 585) out = -7;
	 	 	 else if (in >= 586 && in <= 682) out = -6;
	 	 	 else if (in >= 683 && in <= 819) out = -5;
	 	 	 else if (in >= 820 && in <= 1024) out = -4;
	 	 	 else if (in >= 1025 && in <= 1365) out = -3;
	 	 	 else if (in >= 1366 && in <= 2048) out = -2;
	 	 	 else if (in >= 2049 && in <= 4095) out = -1;
	 	 	else out=0;
	 endmodule
